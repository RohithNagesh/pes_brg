magic
tech sky130A
magscale 1 2
timestamp 1699008247
<< viali >>
rect 6469 10217 6503 10251
rect 5457 10149 5491 10183
rect 7665 10149 7699 10183
rect 2513 10013 2547 10047
rect 2789 10013 2823 10047
rect 4353 10013 4387 10047
rect 4537 10013 4571 10047
rect 5181 10013 5215 10047
rect 5457 10013 5491 10047
rect 7573 10013 7607 10047
rect 7665 10013 7699 10047
rect 7941 10013 7975 10047
rect 8217 10013 8251 10047
rect 6745 9945 6779 9979
rect 7297 9945 7331 9979
rect 7481 9945 7515 9979
rect 2513 9877 2547 9911
rect 3801 9877 3835 9911
rect 4629 9877 4663 9911
rect 5273 9877 5307 9911
rect 7573 9877 7607 9911
rect 7849 9877 7883 9911
rect 8125 9877 8159 9911
rect 1593 9673 1627 9707
rect 6193 9673 6227 9707
rect 7656 9605 7690 9639
rect 1409 9537 1443 9571
rect 1501 9537 1535 9571
rect 2136 9537 2170 9571
rect 3341 9537 3375 9571
rect 3608 9537 3642 9571
rect 4813 9537 4847 9571
rect 5080 9537 5114 9571
rect 7113 9537 7147 9571
rect 7205 9537 7239 9571
rect 7389 9537 7423 9571
rect 1777 9469 1811 9503
rect 1869 9469 1903 9503
rect 7021 9469 7055 9503
rect 1501 9333 1535 9367
rect 3249 9333 3283 9367
rect 4721 9333 4755 9367
rect 6377 9333 6411 9367
rect 8769 9333 8803 9367
rect 2881 9129 2915 9163
rect 6561 9129 6595 9163
rect 6653 9129 6687 9163
rect 7113 9129 7147 9163
rect 7297 9129 7331 9163
rect 7389 9129 7423 9163
rect 4905 9061 4939 9095
rect 5549 9061 5583 9095
rect 5825 9061 5859 9095
rect 5457 8993 5491 9027
rect 6745 8993 6779 9027
rect 7205 8993 7239 9027
rect 1409 8925 1443 8959
rect 3065 8925 3099 8959
rect 3157 8925 3191 8959
rect 3249 8925 3283 8959
rect 3525 8925 3559 8959
rect 4077 8925 4111 8959
rect 4169 8925 4203 8959
rect 4261 8925 4295 8959
rect 4445 8925 4479 8959
rect 5181 8925 5215 8959
rect 5641 8925 5675 8959
rect 5733 8925 5767 8959
rect 6101 8925 6135 8959
rect 6469 8925 6503 8959
rect 6837 8925 6871 8959
rect 7665 8925 7699 8959
rect 8585 8925 8619 8959
rect 1654 8857 1688 8891
rect 3387 8857 3421 8891
rect 4537 8857 4571 8891
rect 4721 8857 4755 8891
rect 5387 8857 5421 8891
rect 7389 8857 7423 8891
rect 8033 8857 8067 8891
rect 2789 8789 2823 8823
rect 3801 8789 3835 8823
rect 5273 8789 5307 8823
rect 5825 8789 5859 8823
rect 5917 8789 5951 8823
rect 6929 8789 6963 8823
rect 7573 8789 7607 8823
rect 1409 8585 1443 8619
rect 2881 8585 2915 8619
rect 3249 8585 3283 8619
rect 4353 8585 4387 8619
rect 5733 8585 5767 8619
rect 6469 8585 6503 8619
rect 7205 8585 7239 8619
rect 8953 8585 8987 8619
rect 1685 8517 1719 8551
rect 6837 8517 6871 8551
rect 7021 8517 7055 8551
rect 7818 8517 7852 8551
rect 1593 8449 1627 8483
rect 1777 8449 1811 8483
rect 1915 8449 1949 8483
rect 2145 8449 2179 8483
rect 3801 8449 3835 8483
rect 4077 8449 4111 8483
rect 4169 8449 4203 8483
rect 4445 8449 4479 8483
rect 6377 8449 6411 8483
rect 6653 8449 6687 8483
rect 6929 8449 6963 8483
rect 7297 8449 7331 8483
rect 7481 8449 7515 8483
rect 2053 8381 2087 8415
rect 2789 8381 2823 8415
rect 3065 8381 3099 8415
rect 3157 8381 3191 8415
rect 3433 8381 3467 8415
rect 3525 8381 3559 8415
rect 7573 8381 7607 8415
rect 3893 8245 3927 8279
rect 1777 8041 1811 8075
rect 3617 8041 3651 8075
rect 5365 8041 5399 8075
rect 5733 8041 5767 8075
rect 7205 8041 7239 8075
rect 7297 8041 7331 8075
rect 7481 8041 7515 8075
rect 7757 8041 7791 8075
rect 3801 7973 3835 8007
rect 3065 7905 3099 7939
rect 4721 7905 4755 7939
rect 5089 7905 5123 7939
rect 2237 7837 2271 7871
rect 2421 7837 2455 7871
rect 2697 7837 2731 7871
rect 3341 7837 3375 7871
rect 3985 7837 4019 7871
rect 5181 7837 5215 7871
rect 5641 7837 5675 7871
rect 5825 7837 5859 7871
rect 6101 7837 6135 7871
rect 6285 7837 6319 7871
rect 6653 7837 6687 7871
rect 6745 7837 6779 7871
rect 6837 7837 6871 7871
rect 7021 7837 7055 7871
rect 7481 7837 7515 7871
rect 7665 7837 7699 7871
rect 7757 7837 7791 7871
rect 7849 7837 7883 7871
rect 8309 7837 8343 7871
rect 1593 7769 1627 7803
rect 2605 7769 2639 7803
rect 3249 7769 3283 7803
rect 8033 7769 8067 7803
rect 1793 7701 1827 7735
rect 1961 7701 1995 7735
rect 3433 7701 3467 7735
rect 8217 7701 8251 7735
rect 5365 7497 5399 7531
rect 6561 7497 6595 7531
rect 7021 7497 7055 7531
rect 8217 7497 8251 7531
rect 6101 7429 6135 7463
rect 1409 7361 1443 7395
rect 1676 7361 1710 7395
rect 3617 7361 3651 7395
rect 4261 7361 4295 7395
rect 4353 7361 4387 7395
rect 5089 7361 5123 7395
rect 5365 7361 5399 7395
rect 5457 7361 5491 7395
rect 5641 7361 5675 7395
rect 5733 7361 5767 7395
rect 5825 7361 5859 7395
rect 6009 7361 6043 7395
rect 6193 7361 6227 7395
rect 6377 7361 6411 7395
rect 6745 7361 6779 7395
rect 7297 7361 7331 7395
rect 7389 7361 7423 7395
rect 2973 7293 3007 7327
rect 3157 7293 3191 7327
rect 3249 7293 3283 7327
rect 3341 7293 3375 7327
rect 3433 7293 3467 7327
rect 7021 7293 7055 7327
rect 7113 7293 7147 7327
rect 8033 7293 8067 7327
rect 8769 7293 8803 7327
rect 2789 7225 2823 7259
rect 4997 7225 5031 7259
rect 7205 7225 7239 7259
rect 6837 7157 6871 7191
rect 7481 7157 7515 7191
rect 1777 6953 1811 6987
rect 2697 6953 2731 6987
rect 8769 6953 8803 6987
rect 1409 6885 1443 6919
rect 2881 6885 2915 6919
rect 5457 6885 5491 6919
rect 1961 6817 1995 6851
rect 7389 6817 7423 6851
rect 1593 6749 1627 6783
rect 1685 6749 1719 6783
rect 2053 6749 2087 6783
rect 2329 6749 2363 6783
rect 3249 6749 3283 6783
rect 3801 6749 3835 6783
rect 3893 6749 3927 6783
rect 4077 6749 4111 6783
rect 4261 6749 4295 6783
rect 4537 6749 4571 6783
rect 4905 6749 4939 6783
rect 5089 6749 5123 6783
rect 5365 6749 5399 6783
rect 5733 6749 5767 6783
rect 6101 6749 6135 6783
rect 7021 6749 7055 6783
rect 7205 6749 7239 6783
rect 7297 6749 7331 6783
rect 7656 6749 7690 6783
rect 1409 6681 1443 6715
rect 2421 6681 2455 6715
rect 2605 6681 2639 6715
rect 4997 6681 5031 6715
rect 6377 6681 6411 6715
rect 6561 6681 6595 6715
rect 3341 6613 3375 6647
rect 6745 6613 6779 6647
rect 6837 6613 6871 6647
rect 2145 6409 2179 6443
rect 2605 6409 2639 6443
rect 3249 6409 3283 6443
rect 5733 6409 5767 6443
rect 6929 6409 6963 6443
rect 8861 6409 8895 6443
rect 1409 6341 1443 6375
rect 4445 6341 4479 6375
rect 7726 6341 7760 6375
rect 1639 6307 1673 6341
rect 2237 6273 2271 6307
rect 3065 6273 3099 6307
rect 3341 6273 3375 6307
rect 3893 6273 3927 6307
rect 4169 6273 4203 6307
rect 6469 6273 6503 6307
rect 6561 6273 6595 6307
rect 6653 6273 6687 6307
rect 6745 6273 6779 6307
rect 7113 6273 7147 6307
rect 7205 6273 7239 6307
rect 7389 6273 7423 6307
rect 7481 6273 7515 6307
rect 1961 6205 1995 6239
rect 2789 6205 2823 6239
rect 2973 6205 3007 6239
rect 3433 6205 3467 6239
rect 3525 6205 3559 6239
rect 3709 6205 3743 6239
rect 3801 6205 3835 6239
rect 3985 6205 4019 6239
rect 1777 6137 1811 6171
rect 4353 6137 4387 6171
rect 1593 6069 1627 6103
rect 7297 6069 7331 6103
rect 3157 5865 3191 5899
rect 5181 5865 5215 5899
rect 5365 5865 5399 5899
rect 6469 5865 6503 5899
rect 7481 5865 7515 5899
rect 2789 5797 2823 5831
rect 4997 5797 5031 5831
rect 3525 5729 3559 5763
rect 4353 5729 4387 5763
rect 4721 5729 4755 5763
rect 5641 5729 5675 5763
rect 5733 5729 5767 5763
rect 5825 5729 5859 5763
rect 7757 5729 7791 5763
rect 1409 5661 1443 5695
rect 1676 5661 1710 5695
rect 2881 5661 2915 5695
rect 3341 5661 3375 5695
rect 3617 5661 3651 5695
rect 4077 5661 4111 5695
rect 4261 5661 4295 5695
rect 4629 5661 4663 5695
rect 5457 5661 5491 5695
rect 5917 5661 5951 5695
rect 6377 5661 6411 5695
rect 6653 5661 6687 5695
rect 6929 5661 6963 5695
rect 7021 5661 7055 5695
rect 7389 5661 7423 5695
rect 8125 5661 8159 5695
rect 8401 5661 8435 5695
rect 8677 5661 8711 5695
rect 4537 5593 4571 5627
rect 7640 5593 7674 5627
rect 8217 5593 8251 5627
rect 8585 5593 8619 5627
rect 2973 5525 3007 5559
rect 6101 5525 6135 5559
rect 7849 5525 7883 5559
rect 3157 5321 3191 5355
rect 7941 5321 7975 5355
rect 8033 5321 8067 5355
rect 8217 5321 8251 5355
rect 8677 5321 8711 5355
rect 1409 5185 1443 5219
rect 1676 5185 1710 5219
rect 2973 5185 3007 5219
rect 3157 5185 3191 5219
rect 3893 5185 3927 5219
rect 4353 5185 4387 5219
rect 4629 5185 4663 5219
rect 4905 5185 4939 5219
rect 4997 5185 5031 5219
rect 5733 5185 5767 5219
rect 5917 5185 5951 5219
rect 6377 5185 6411 5219
rect 6561 5185 6595 5219
rect 6837 5185 6871 5219
rect 7113 5185 7147 5219
rect 7297 5185 7331 5219
rect 7757 5185 7791 5219
rect 8125 5185 8159 5219
rect 8217 5185 8251 5219
rect 8585 5185 8619 5219
rect 8769 5185 8803 5219
rect 3617 5117 3651 5151
rect 8309 5117 8343 5151
rect 8493 5117 8527 5151
rect 2789 4981 2823 5015
rect 6469 4981 6503 5015
rect 7481 4981 7515 5015
rect 7849 4981 7883 5015
rect 1685 4777 1719 4811
rect 2789 4777 2823 4811
rect 6193 4777 6227 4811
rect 5549 4709 5583 4743
rect 3157 4641 3191 4675
rect 3985 4641 4019 4675
rect 5089 4641 5123 4675
rect 5181 4641 5215 4675
rect 5365 4641 5399 4675
rect 5641 4641 5675 4675
rect 1869 4573 1903 4607
rect 2145 4573 2179 4607
rect 2329 4573 2363 4607
rect 2513 4573 2547 4607
rect 2605 4573 2639 4607
rect 3571 4573 3605 4607
rect 3893 4573 3927 4607
rect 4077 4573 4111 4607
rect 4261 4573 4295 4607
rect 4629 4573 4663 4607
rect 4997 4573 5031 4607
rect 5825 4573 5859 4607
rect 5917 4573 5951 4607
rect 6009 4573 6043 4607
rect 6653 4573 6687 4607
rect 7113 4573 7147 4607
rect 7205 4573 7239 4607
rect 7297 4573 7331 4607
rect 7389 4573 7423 4607
rect 7573 4573 7607 4607
rect 8033 4573 8067 4607
rect 8217 4573 8251 4607
rect 8493 4573 8527 4607
rect 5273 4505 5307 4539
rect 6469 4505 6503 4539
rect 7849 4505 7883 4539
rect 1961 4437 1995 4471
rect 4261 4437 4295 4471
rect 6285 4437 6319 4471
rect 6929 4437 6963 4471
rect 6101 4233 6135 4267
rect 7941 4233 7975 4267
rect 5457 4165 5491 4199
rect 1409 4097 1443 4131
rect 1676 4097 1710 4131
rect 5641 4097 5675 4131
rect 5825 4097 5859 4131
rect 6193 4097 6227 4131
rect 7113 4097 7147 4131
rect 7573 4097 7607 4131
rect 8401 4097 8435 4131
rect 3433 4029 3467 4063
rect 6837 4029 6871 4063
rect 8125 4029 8159 4063
rect 8217 4029 8251 4063
rect 8309 4029 8343 4063
rect 4169 3961 4203 3995
rect 6561 3961 6595 3995
rect 2789 3893 2823 3927
rect 2881 3893 2915 3927
rect 5825 3893 5859 3927
rect 6837 3893 6871 3927
rect 7297 3893 7331 3927
rect 1593 3689 1627 3723
rect 2053 3689 2087 3723
rect 2145 3689 2179 3723
rect 6377 3689 6411 3723
rect 7021 3689 7055 3723
rect 8125 3689 8159 3723
rect 3985 3621 4019 3655
rect 4169 3621 4203 3655
rect 4629 3621 4663 3655
rect 6469 3621 6503 3655
rect 8309 3621 8343 3655
rect 1961 3553 1995 3587
rect 3893 3553 3927 3587
rect 4905 3553 4939 3587
rect 7665 3553 7699 3587
rect 1409 3485 1443 3519
rect 2237 3485 2271 3519
rect 2513 3485 2547 3519
rect 2697 3485 2731 3519
rect 3341 3485 3375 3519
rect 4169 3485 4203 3519
rect 4353 3485 4387 3519
rect 4537 3485 4571 3519
rect 4813 3485 4847 3519
rect 4997 3485 5031 3519
rect 5181 3485 5215 3519
rect 5457 3485 5491 3519
rect 5641 3485 5675 3519
rect 5917 3485 5951 3519
rect 6285 3485 6319 3519
rect 6745 3485 6779 3519
rect 6837 3485 6871 3519
rect 7941 3485 7975 3519
rect 8033 3485 8067 3519
rect 8217 3485 8251 3519
rect 8309 3485 8343 3519
rect 8493 3485 8527 3519
rect 4261 3417 4295 3451
rect 5273 3417 5307 3451
rect 2329 3349 2363 3383
rect 2789 3349 2823 3383
rect 5089 3349 5123 3383
rect 7849 3349 7883 3383
rect 4077 3145 4111 3179
rect 4169 3145 4203 3179
rect 4445 3145 4479 3179
rect 7941 3145 7975 3179
rect 3801 3077 3835 3111
rect 3893 3077 3927 3111
rect 6622 3077 6656 3111
rect 1593 3009 1627 3043
rect 1860 3009 1894 3043
rect 3157 3009 3191 3043
rect 3249 3009 3283 3043
rect 3617 3009 3651 3043
rect 4261 3009 4295 3043
rect 5742 3009 5776 3043
rect 6009 3009 6043 3043
rect 6377 3009 6411 3043
rect 8493 2941 8527 2975
rect 7757 2873 7791 2907
rect 2973 2805 3007 2839
rect 4629 2805 4663 2839
rect 1777 2601 1811 2635
rect 2145 2601 2179 2635
rect 2421 2601 2455 2635
rect 3341 2601 3375 2635
rect 3985 2601 4019 2635
rect 4445 2601 4479 2635
rect 5733 2601 5767 2635
rect 6193 2601 6227 2635
rect 8033 2601 8067 2635
rect 2697 2533 2731 2567
rect 5825 2533 5859 2567
rect 1869 2465 1903 2499
rect 3157 2465 3191 2499
rect 4077 2465 4111 2499
rect 6653 2465 6687 2499
rect 1593 2397 1627 2431
rect 1685 2397 1719 2431
rect 2053 2397 2087 2431
rect 2513 2397 2547 2431
rect 2789 2397 2823 2431
rect 3065 2397 3099 2431
rect 3249 2397 3283 2431
rect 3525 2397 3559 2431
rect 3801 2397 3835 2431
rect 3985 2397 4019 2431
rect 4261 2397 4295 2431
rect 4721 2397 4755 2431
rect 5273 2397 5307 2431
rect 5365 2397 5399 2431
rect 5457 2397 5491 2431
rect 5917 2397 5951 2431
rect 6009 2397 6043 2431
rect 6920 2397 6954 2431
<< metal1 >>
rect 1104 10362 9292 10384
rect 1104 10310 1973 10362
rect 2025 10310 2037 10362
rect 2089 10310 2101 10362
rect 2153 10310 2165 10362
rect 2217 10310 2229 10362
rect 2281 10310 4020 10362
rect 4072 10310 4084 10362
rect 4136 10310 4148 10362
rect 4200 10310 4212 10362
rect 4264 10310 4276 10362
rect 4328 10310 6067 10362
rect 6119 10310 6131 10362
rect 6183 10310 6195 10362
rect 6247 10310 6259 10362
rect 6311 10310 6323 10362
rect 6375 10310 8114 10362
rect 8166 10310 8178 10362
rect 8230 10310 8242 10362
rect 8294 10310 8306 10362
rect 8358 10310 8370 10362
rect 8422 10310 9292 10362
rect 1104 10288 9292 10310
rect 5810 10208 5816 10260
rect 5868 10248 5874 10260
rect 6457 10251 6515 10257
rect 6457 10248 6469 10251
rect 5868 10220 6469 10248
rect 5868 10208 5874 10220
rect 6457 10217 6469 10220
rect 6503 10217 6515 10251
rect 6457 10211 6515 10217
rect 5350 10140 5356 10192
rect 5408 10180 5414 10192
rect 5445 10183 5503 10189
rect 5445 10180 5457 10183
rect 5408 10152 5457 10180
rect 5408 10140 5414 10152
rect 5445 10149 5457 10152
rect 5491 10149 5503 10183
rect 5445 10143 5503 10149
rect 7650 10140 7656 10192
rect 7708 10140 7714 10192
rect 7282 10072 7288 10124
rect 7340 10112 7346 10124
rect 7340 10084 7696 10112
rect 7340 10072 7346 10084
rect 2038 10004 2044 10056
rect 2096 10044 2102 10056
rect 2501 10047 2559 10053
rect 2501 10044 2513 10047
rect 2096 10016 2513 10044
rect 2096 10004 2102 10016
rect 2501 10013 2513 10016
rect 2547 10013 2559 10047
rect 2501 10007 2559 10013
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10044 2835 10047
rect 2958 10044 2964 10056
rect 2823 10016 2964 10044
rect 2823 10013 2835 10016
rect 2777 10007 2835 10013
rect 2958 10004 2964 10016
rect 3016 10004 3022 10056
rect 3234 10004 3240 10056
rect 3292 10044 3298 10056
rect 4341 10047 4399 10053
rect 4341 10044 4353 10047
rect 3292 10016 4353 10044
rect 3292 10004 3298 10016
rect 4341 10013 4353 10016
rect 4387 10044 4399 10047
rect 4525 10047 4583 10053
rect 4525 10044 4537 10047
rect 4387 10016 4537 10044
rect 4387 10013 4399 10016
rect 4341 10007 4399 10013
rect 4525 10013 4537 10016
rect 4571 10013 4583 10047
rect 4525 10007 4583 10013
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10044 5227 10047
rect 5258 10044 5264 10056
rect 5215 10016 5264 10044
rect 5215 10013 5227 10016
rect 5169 10007 5227 10013
rect 5258 10004 5264 10016
rect 5316 10004 5322 10056
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10044 5503 10047
rect 7190 10044 7196 10056
rect 5491 10016 7196 10044
rect 5491 10013 5503 10016
rect 5445 10007 5503 10013
rect 7190 10004 7196 10016
rect 7248 10004 7254 10056
rect 7558 10004 7564 10056
rect 7616 10004 7622 10056
rect 7668 10053 7696 10084
rect 7653 10047 7711 10053
rect 7653 10013 7665 10047
rect 7699 10013 7711 10047
rect 7929 10047 7987 10053
rect 7929 10044 7941 10047
rect 7653 10007 7711 10013
rect 7760 10016 7941 10044
rect 6178 9936 6184 9988
rect 6236 9976 6242 9988
rect 6733 9979 6791 9985
rect 6733 9976 6745 9979
rect 6236 9948 6745 9976
rect 6236 9936 6242 9948
rect 6733 9945 6745 9948
rect 6779 9945 6791 9979
rect 6733 9939 6791 9945
rect 7098 9936 7104 9988
rect 7156 9976 7162 9988
rect 7285 9979 7343 9985
rect 7285 9976 7297 9979
rect 7156 9948 7297 9976
rect 7156 9936 7162 9948
rect 7285 9945 7297 9948
rect 7331 9945 7343 9979
rect 7285 9939 7343 9945
rect 7466 9936 7472 9988
rect 7524 9936 7530 9988
rect 2498 9868 2504 9920
rect 2556 9868 2562 9920
rect 3418 9868 3424 9920
rect 3476 9908 3482 9920
rect 3789 9911 3847 9917
rect 3789 9908 3801 9911
rect 3476 9880 3801 9908
rect 3476 9868 3482 9880
rect 3789 9877 3801 9880
rect 3835 9877 3847 9911
rect 3789 9871 3847 9877
rect 4522 9868 4528 9920
rect 4580 9908 4586 9920
rect 4617 9911 4675 9917
rect 4617 9908 4629 9911
rect 4580 9880 4629 9908
rect 4580 9868 4586 9880
rect 4617 9877 4629 9880
rect 4663 9877 4675 9911
rect 4617 9871 4675 9877
rect 5074 9868 5080 9920
rect 5132 9908 5138 9920
rect 5261 9911 5319 9917
rect 5261 9908 5273 9911
rect 5132 9880 5273 9908
rect 5132 9868 5138 9880
rect 5261 9877 5273 9880
rect 5307 9877 5319 9911
rect 5261 9871 5319 9877
rect 7561 9911 7619 9917
rect 7561 9877 7573 9911
rect 7607 9908 7619 9911
rect 7760 9908 7788 10016
rect 7929 10013 7941 10016
rect 7975 10013 7987 10047
rect 7929 10007 7987 10013
rect 8205 10047 8263 10053
rect 8205 10013 8217 10047
rect 8251 10013 8263 10047
rect 8205 10007 8263 10013
rect 8018 9936 8024 9988
rect 8076 9976 8082 9988
rect 8220 9976 8248 10007
rect 8076 9948 8248 9976
rect 8076 9936 8082 9948
rect 7607 9880 7788 9908
rect 7607 9877 7619 9880
rect 7561 9871 7619 9877
rect 7834 9868 7840 9920
rect 7892 9908 7898 9920
rect 8113 9911 8171 9917
rect 8113 9908 8125 9911
rect 7892 9880 8125 9908
rect 7892 9868 7898 9880
rect 8113 9877 8125 9880
rect 8159 9877 8171 9911
rect 8113 9871 8171 9877
rect 1104 9818 9292 9840
rect 1104 9766 2633 9818
rect 2685 9766 2697 9818
rect 2749 9766 2761 9818
rect 2813 9766 2825 9818
rect 2877 9766 2889 9818
rect 2941 9766 4680 9818
rect 4732 9766 4744 9818
rect 4796 9766 4808 9818
rect 4860 9766 4872 9818
rect 4924 9766 4936 9818
rect 4988 9766 6727 9818
rect 6779 9766 6791 9818
rect 6843 9766 6855 9818
rect 6907 9766 6919 9818
rect 6971 9766 6983 9818
rect 7035 9766 8774 9818
rect 8826 9766 8838 9818
rect 8890 9766 8902 9818
rect 8954 9766 8966 9818
rect 9018 9766 9030 9818
rect 9082 9766 9292 9818
rect 1104 9744 9292 9766
rect 1578 9664 1584 9716
rect 1636 9664 1642 9716
rect 2038 9704 2044 9716
rect 1688 9676 2044 9704
rect 1688 9648 1716 9676
rect 2038 9664 2044 9676
rect 2096 9664 2102 9716
rect 6178 9664 6184 9716
rect 6236 9664 6242 9716
rect 1670 9636 1676 9648
rect 1412 9608 1676 9636
rect 1412 9577 1440 9608
rect 1670 9596 1676 9608
rect 1728 9596 1734 9648
rect 5718 9636 5724 9648
rect 1872 9608 5724 9636
rect 1397 9571 1455 9577
rect 1397 9537 1409 9571
rect 1443 9537 1455 9571
rect 1397 9531 1455 9537
rect 1489 9571 1547 9577
rect 1489 9537 1501 9571
rect 1535 9537 1547 9571
rect 1489 9531 1547 9537
rect 1504 9500 1532 9531
rect 1578 9528 1584 9580
rect 1636 9568 1642 9580
rect 1872 9568 1900 9608
rect 1636 9540 1900 9568
rect 1636 9528 1642 9540
rect 1504 9472 1716 9500
rect 1489 9367 1547 9373
rect 1489 9333 1501 9367
rect 1535 9364 1547 9367
rect 1578 9364 1584 9376
rect 1535 9336 1584 9364
rect 1535 9333 1547 9336
rect 1489 9327 1547 9333
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 1688 9364 1716 9472
rect 1762 9460 1768 9512
rect 1820 9460 1826 9512
rect 1872 9509 1900 9540
rect 2124 9571 2182 9577
rect 2124 9537 2136 9571
rect 2170 9568 2182 9571
rect 2866 9568 2872 9580
rect 2170 9540 2872 9568
rect 2170 9537 2182 9540
rect 2124 9531 2182 9537
rect 2866 9528 2872 9540
rect 2924 9528 2930 9580
rect 3344 9577 3372 9608
rect 3329 9571 3387 9577
rect 3329 9537 3341 9571
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 3596 9571 3654 9577
rect 3596 9537 3608 9571
rect 3642 9568 3654 9571
rect 4338 9568 4344 9580
rect 3642 9540 4344 9568
rect 3642 9537 3654 9540
rect 3596 9531 3654 9537
rect 4338 9528 4344 9540
rect 4396 9528 4402 9580
rect 4816 9577 4844 9608
rect 5718 9596 5724 9608
rect 5776 9636 5782 9648
rect 7650 9645 7656 9648
rect 7644 9636 7656 9645
rect 5776 9608 7420 9636
rect 7611 9608 7656 9636
rect 5776 9596 5782 9608
rect 7392 9580 7420 9608
rect 7644 9599 7656 9608
rect 7650 9596 7656 9599
rect 7708 9596 7714 9648
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 5068 9571 5126 9577
rect 5068 9537 5080 9571
rect 5114 9568 5126 9571
rect 5442 9568 5448 9580
rect 5114 9540 5448 9568
rect 5114 9537 5126 9540
rect 5068 9531 5126 9537
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 6178 9528 6184 9580
rect 6236 9568 6242 9580
rect 7101 9571 7159 9577
rect 7101 9568 7113 9571
rect 6236 9540 7113 9568
rect 6236 9528 6242 9540
rect 7101 9537 7113 9540
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 7190 9528 7196 9580
rect 7248 9528 7254 9580
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9469 1915 9503
rect 1857 9463 1915 9469
rect 7009 9503 7067 9509
rect 7009 9469 7021 9503
rect 7055 9500 7067 9503
rect 7208 9500 7236 9528
rect 7055 9472 7236 9500
rect 7055 9469 7067 9472
rect 7009 9463 7067 9469
rect 2958 9364 2964 9376
rect 1688 9336 2964 9364
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 3234 9324 3240 9376
rect 3292 9324 3298 9376
rect 4522 9324 4528 9376
rect 4580 9364 4586 9376
rect 4709 9367 4767 9373
rect 4709 9364 4721 9367
rect 4580 9336 4721 9364
rect 4580 9324 4586 9336
rect 4709 9333 4721 9336
rect 4755 9333 4767 9367
rect 4709 9327 4767 9333
rect 5534 9324 5540 9376
rect 5592 9364 5598 9376
rect 6365 9367 6423 9373
rect 6365 9364 6377 9367
rect 5592 9336 6377 9364
rect 5592 9324 5598 9336
rect 6365 9333 6377 9336
rect 6411 9333 6423 9367
rect 6365 9327 6423 9333
rect 8018 9324 8024 9376
rect 8076 9364 8082 9376
rect 8757 9367 8815 9373
rect 8757 9364 8769 9367
rect 8076 9336 8769 9364
rect 8076 9324 8082 9336
rect 8757 9333 8769 9336
rect 8803 9333 8815 9367
rect 8757 9327 8815 9333
rect 1104 9274 9292 9296
rect 1104 9222 1973 9274
rect 2025 9222 2037 9274
rect 2089 9222 2101 9274
rect 2153 9222 2165 9274
rect 2217 9222 2229 9274
rect 2281 9222 4020 9274
rect 4072 9222 4084 9274
rect 4136 9222 4148 9274
rect 4200 9222 4212 9274
rect 4264 9222 4276 9274
rect 4328 9222 6067 9274
rect 6119 9222 6131 9274
rect 6183 9222 6195 9274
rect 6247 9222 6259 9274
rect 6311 9222 6323 9274
rect 6375 9222 8114 9274
rect 8166 9222 8178 9274
rect 8230 9222 8242 9274
rect 8294 9222 8306 9274
rect 8358 9222 8370 9274
rect 8422 9222 9292 9274
rect 1104 9200 9292 9222
rect 2866 9120 2872 9172
rect 2924 9120 2930 9172
rect 5442 9120 5448 9172
rect 5500 9120 5506 9172
rect 5994 9120 6000 9172
rect 6052 9160 6058 9172
rect 6549 9163 6607 9169
rect 6549 9160 6561 9163
rect 6052 9132 6561 9160
rect 6052 9120 6058 9132
rect 6549 9129 6561 9132
rect 6595 9129 6607 9163
rect 6549 9123 6607 9129
rect 6641 9163 6699 9169
rect 6641 9129 6653 9163
rect 6687 9160 6699 9163
rect 6914 9160 6920 9172
rect 6687 9132 6920 9160
rect 6687 9129 6699 9132
rect 6641 9123 6699 9129
rect 6914 9120 6920 9132
rect 6972 9160 6978 9172
rect 7101 9163 7159 9169
rect 7101 9160 7113 9163
rect 6972 9132 7113 9160
rect 6972 9120 6978 9132
rect 7101 9129 7113 9132
rect 7147 9129 7159 9163
rect 7101 9123 7159 9129
rect 7282 9120 7288 9172
rect 7340 9120 7346 9172
rect 7377 9163 7435 9169
rect 7377 9129 7389 9163
rect 7423 9160 7435 9163
rect 7466 9160 7472 9172
rect 7423 9132 7472 9160
rect 7423 9129 7435 9132
rect 7377 9123 7435 9129
rect 7466 9120 7472 9132
rect 7524 9120 7530 9172
rect 3142 9052 3148 9104
rect 3200 9092 3206 9104
rect 4893 9095 4951 9101
rect 4893 9092 4905 9095
rect 3200 9064 4905 9092
rect 3200 9052 3206 9064
rect 4893 9061 4905 9064
rect 4939 9061 4951 9095
rect 5460 9092 5488 9120
rect 5537 9095 5595 9101
rect 5537 9092 5549 9095
rect 5460 9064 5549 9092
rect 4893 9055 4951 9061
rect 5537 9061 5549 9064
rect 5583 9061 5595 9095
rect 5813 9095 5871 9101
rect 5813 9092 5825 9095
rect 5537 9055 5595 9061
rect 5644 9064 5825 9092
rect 5074 9024 5080 9036
rect 3252 8996 5080 9024
rect 1394 8916 1400 8968
rect 1452 8916 1458 8968
rect 3050 8916 3056 8968
rect 3108 8916 3114 8968
rect 3142 8916 3148 8968
rect 3200 8916 3206 8968
rect 3252 8965 3280 8996
rect 3237 8959 3295 8965
rect 3237 8925 3249 8959
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8925 3571 8959
rect 3513 8919 3571 8925
rect 1486 8848 1492 8900
rect 1544 8888 1550 8900
rect 3418 8897 3424 8900
rect 1642 8891 1700 8897
rect 1642 8888 1654 8891
rect 1544 8860 1654 8888
rect 1544 8848 1550 8860
rect 1642 8857 1654 8860
rect 1688 8857 1700 8891
rect 1642 8851 1700 8857
rect 3375 8891 3424 8897
rect 3375 8857 3387 8891
rect 3421 8857 3424 8891
rect 3375 8851 3424 8857
rect 3418 8848 3424 8851
rect 3476 8848 3482 8900
rect 2777 8823 2835 8829
rect 2777 8789 2789 8823
rect 2823 8820 2835 8823
rect 2958 8820 2964 8832
rect 2823 8792 2964 8820
rect 2823 8789 2835 8792
rect 2777 8783 2835 8789
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 3142 8780 3148 8832
rect 3200 8820 3206 8832
rect 3528 8820 3556 8919
rect 3620 8900 3648 8996
rect 3878 8916 3884 8968
rect 3936 8956 3942 8968
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 3936 8928 4077 8956
rect 3936 8916 3942 8928
rect 4065 8925 4077 8928
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 3602 8848 3608 8900
rect 3660 8848 3666 8900
rect 3200 8792 3556 8820
rect 3200 8780 3206 8792
rect 3786 8780 3792 8832
rect 3844 8780 3850 8832
rect 4080 8820 4108 8919
rect 4154 8916 4160 8968
rect 4212 8916 4218 8968
rect 4246 8916 4252 8968
rect 4304 8916 4310 8968
rect 4448 8965 4476 8996
rect 5074 8984 5080 8996
rect 5132 9024 5138 9036
rect 5445 9027 5503 9033
rect 5132 8996 5304 9024
rect 5132 8984 5138 8996
rect 4433 8959 4491 8965
rect 4433 8925 4445 8959
rect 4479 8925 4491 8959
rect 4433 8919 4491 8925
rect 5166 8916 5172 8968
rect 5224 8916 5230 8968
rect 5276 8956 5304 8996
rect 5445 8993 5457 9027
rect 5491 9024 5503 9027
rect 5644 9024 5672 9064
rect 5813 9061 5825 9064
rect 5859 9061 5871 9095
rect 5813 9055 5871 9061
rect 6472 9064 7144 9092
rect 5491 8996 5672 9024
rect 5491 8993 5503 8996
rect 5445 8987 5503 8993
rect 5276 8928 5598 8956
rect 4172 8888 4200 8916
rect 5570 8900 5598 8928
rect 5626 8916 5632 8968
rect 5684 8916 5690 8968
rect 5721 8959 5779 8965
rect 5721 8925 5733 8959
rect 5767 8925 5779 8959
rect 5721 8922 5779 8925
rect 6089 8959 6147 8965
rect 6089 8925 6101 8959
rect 6135 8956 6147 8959
rect 6178 8956 6184 8968
rect 6135 8928 6184 8956
rect 6135 8925 6147 8928
rect 5721 8919 5856 8922
rect 6089 8919 6147 8925
rect 4525 8891 4583 8897
rect 4525 8888 4537 8891
rect 4172 8860 4537 8888
rect 4525 8857 4537 8860
rect 4571 8857 4583 8891
rect 4525 8851 4583 8857
rect 4709 8891 4767 8897
rect 4709 8857 4721 8891
rect 4755 8857 4767 8891
rect 4709 8851 4767 8857
rect 4614 8820 4620 8832
rect 4080 8792 4620 8820
rect 4614 8780 4620 8792
rect 4672 8820 4678 8832
rect 4724 8820 4752 8851
rect 5350 8848 5356 8900
rect 5408 8897 5414 8900
rect 5408 8891 5433 8897
rect 5421 8857 5433 8891
rect 5408 8851 5433 8857
rect 5408 8848 5414 8851
rect 5534 8848 5540 8900
rect 5592 8888 5598 8900
rect 5745 8894 5856 8919
rect 6178 8916 6184 8928
rect 6236 8916 6242 8968
rect 6270 8916 6276 8968
rect 6328 8956 6334 8968
rect 6472 8965 6500 9064
rect 6733 9027 6791 9033
rect 6733 9024 6745 9027
rect 6656 8996 6745 9024
rect 6656 8968 6684 8996
rect 6733 8993 6745 8996
rect 6779 8993 6791 9027
rect 6733 8987 6791 8993
rect 6457 8959 6515 8965
rect 6457 8956 6469 8959
rect 6328 8928 6469 8956
rect 6328 8916 6334 8928
rect 6457 8925 6469 8928
rect 6503 8925 6515 8959
rect 6457 8919 6515 8925
rect 6638 8916 6644 8968
rect 6696 8916 6702 8968
rect 6822 8916 6828 8968
rect 6880 8916 6886 8968
rect 5745 8888 5773 8894
rect 5592 8860 5773 8888
rect 5828 8888 5856 8894
rect 7116 8888 7144 9064
rect 7193 9027 7251 9033
rect 7193 8993 7205 9027
rect 7239 9024 7251 9027
rect 7834 9024 7840 9036
rect 7239 8996 7840 9024
rect 7239 8993 7251 8996
rect 7193 8987 7251 8993
rect 7834 8984 7840 8996
rect 7892 8984 7898 9036
rect 7650 8916 7656 8968
rect 7708 8956 7714 8968
rect 8573 8959 8631 8965
rect 8573 8956 8585 8959
rect 7708 8928 8585 8956
rect 7708 8916 7714 8928
rect 8573 8925 8585 8928
rect 8619 8925 8631 8959
rect 8573 8919 8631 8925
rect 7377 8891 7435 8897
rect 7377 8888 7389 8891
rect 5828 8860 6960 8888
rect 7116 8860 7389 8888
rect 5592 8848 5598 8860
rect 4672 8792 4752 8820
rect 5261 8823 5319 8829
rect 4672 8780 4678 8792
rect 5261 8789 5273 8823
rect 5307 8820 5319 8823
rect 5810 8820 5816 8832
rect 5307 8792 5816 8820
rect 5307 8789 5319 8792
rect 5261 8783 5319 8789
rect 5810 8780 5816 8792
rect 5868 8780 5874 8832
rect 5902 8780 5908 8832
rect 5960 8780 5966 8832
rect 6932 8829 6960 8860
rect 7377 8857 7389 8860
rect 7423 8857 7435 8891
rect 8021 8891 8079 8897
rect 8021 8888 8033 8891
rect 7377 8851 7435 8857
rect 7484 8860 8033 8888
rect 6917 8823 6975 8829
rect 6917 8789 6929 8823
rect 6963 8789 6975 8823
rect 6917 8783 6975 8789
rect 7098 8780 7104 8832
rect 7156 8820 7162 8832
rect 7484 8820 7512 8860
rect 8021 8857 8033 8860
rect 8067 8857 8079 8891
rect 8021 8851 8079 8857
rect 7156 8792 7512 8820
rect 7561 8823 7619 8829
rect 7156 8780 7162 8792
rect 7561 8789 7573 8823
rect 7607 8820 7619 8823
rect 7834 8820 7840 8832
rect 7607 8792 7840 8820
rect 7607 8789 7619 8792
rect 7561 8783 7619 8789
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 1104 8730 9292 8752
rect 1104 8678 2633 8730
rect 2685 8678 2697 8730
rect 2749 8678 2761 8730
rect 2813 8678 2825 8730
rect 2877 8678 2889 8730
rect 2941 8678 4680 8730
rect 4732 8678 4744 8730
rect 4796 8678 4808 8730
rect 4860 8678 4872 8730
rect 4924 8678 4936 8730
rect 4988 8678 6727 8730
rect 6779 8678 6791 8730
rect 6843 8678 6855 8730
rect 6907 8678 6919 8730
rect 6971 8678 6983 8730
rect 7035 8678 8774 8730
rect 8826 8678 8838 8730
rect 8890 8678 8902 8730
rect 8954 8678 8966 8730
rect 9018 8678 9030 8730
rect 9082 8678 9292 8730
rect 1104 8656 9292 8678
rect 1397 8619 1455 8625
rect 1397 8585 1409 8619
rect 1443 8616 1455 8619
rect 1486 8616 1492 8628
rect 1443 8588 1492 8616
rect 1443 8585 1455 8588
rect 1397 8579 1455 8585
rect 1486 8576 1492 8588
rect 1544 8576 1550 8628
rect 1578 8576 1584 8628
rect 1636 8576 1642 8628
rect 2869 8619 2927 8625
rect 2869 8585 2881 8619
rect 2915 8616 2927 8619
rect 3050 8616 3056 8628
rect 2915 8588 3056 8616
rect 2915 8585 2927 8588
rect 2869 8579 2927 8585
rect 3050 8576 3056 8588
rect 3108 8576 3114 8628
rect 3237 8619 3295 8625
rect 3237 8585 3249 8619
rect 3283 8585 3295 8619
rect 3237 8579 3295 8585
rect 1596 8548 1624 8576
rect 1673 8551 1731 8557
rect 1673 8548 1685 8551
rect 1596 8520 1685 8548
rect 1673 8517 1685 8520
rect 1719 8517 1731 8551
rect 3142 8548 3148 8560
rect 1673 8511 1731 8517
rect 2424 8520 3148 8548
rect 1302 8440 1308 8492
rect 1360 8480 1366 8492
rect 1581 8483 1639 8489
rect 1581 8480 1593 8483
rect 1360 8452 1593 8480
rect 1360 8440 1366 8452
rect 1581 8449 1593 8452
rect 1627 8449 1639 8483
rect 1581 8443 1639 8449
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8449 1823 8483
rect 1765 8443 1823 8449
rect 1903 8483 1961 8489
rect 1903 8449 1915 8483
rect 1949 8480 1961 8483
rect 2133 8483 2191 8489
rect 2133 8480 2145 8483
rect 1949 8452 2145 8480
rect 1949 8449 1961 8452
rect 1903 8443 1961 8449
rect 2133 8449 2145 8452
rect 2179 8449 2191 8483
rect 2133 8443 2191 8449
rect 1780 8412 1808 8443
rect 2041 8415 2099 8421
rect 1780 8384 1900 8412
rect 1872 8356 1900 8384
rect 2041 8381 2053 8415
rect 2087 8412 2099 8415
rect 2424 8412 2452 8520
rect 3142 8508 3148 8520
rect 3200 8508 3206 8560
rect 3252 8480 3280 8579
rect 3786 8576 3792 8628
rect 3844 8576 3850 8628
rect 4338 8576 4344 8628
rect 4396 8576 4402 8628
rect 5166 8576 5172 8628
rect 5224 8576 5230 8628
rect 5718 8576 5724 8628
rect 5776 8576 5782 8628
rect 6457 8619 6515 8625
rect 6457 8616 6469 8619
rect 6012 8588 6469 8616
rect 3804 8548 3832 8576
rect 5184 8548 5212 8576
rect 5902 8548 5908 8560
rect 3804 8520 4108 8548
rect 5184 8520 5908 8548
rect 2976 8452 3280 8480
rect 2087 8384 2452 8412
rect 2777 8415 2835 8421
rect 2087 8381 2099 8384
rect 2041 8375 2099 8381
rect 2777 8381 2789 8415
rect 2823 8412 2835 8415
rect 2866 8412 2872 8424
rect 2823 8384 2872 8412
rect 2823 8381 2835 8384
rect 2777 8375 2835 8381
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 1854 8304 1860 8356
rect 1912 8304 1918 8356
rect 2976 8288 3004 8452
rect 3326 8440 3332 8492
rect 3384 8480 3390 8492
rect 4080 8489 4108 8520
rect 5902 8508 5908 8520
rect 5960 8508 5966 8560
rect 3789 8483 3847 8489
rect 3789 8480 3801 8483
rect 3384 8452 3801 8480
rect 3384 8440 3390 8452
rect 3789 8449 3801 8452
rect 3835 8449 3847 8483
rect 3789 8443 3847 8449
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8480 4215 8483
rect 4338 8480 4344 8492
rect 4203 8452 4344 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 3053 8415 3111 8421
rect 3053 8381 3065 8415
rect 3099 8381 3111 8415
rect 3053 8375 3111 8381
rect 3145 8415 3203 8421
rect 3145 8381 3157 8415
rect 3191 8412 3203 8415
rect 3191 8384 3372 8412
rect 3191 8381 3203 8384
rect 3145 8375 3203 8381
rect 3068 8344 3096 8375
rect 3234 8344 3240 8356
rect 3068 8316 3240 8344
rect 3234 8304 3240 8316
rect 3292 8304 3298 8356
rect 1486 8236 1492 8288
rect 1544 8276 1550 8288
rect 1946 8276 1952 8288
rect 1544 8248 1952 8276
rect 1544 8236 1550 8248
rect 1946 8236 1952 8248
rect 2004 8276 2010 8288
rect 2958 8276 2964 8288
rect 2004 8248 2964 8276
rect 2004 8236 2010 8248
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 3050 8236 3056 8288
rect 3108 8276 3114 8288
rect 3344 8276 3372 8384
rect 3418 8372 3424 8424
rect 3476 8372 3482 8424
rect 3510 8372 3516 8424
rect 3568 8372 3574 8424
rect 3804 8412 3832 8443
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8480 4491 8483
rect 5442 8480 5448 8492
rect 4479 8452 5448 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 5534 8440 5540 8492
rect 5592 8480 5598 8492
rect 6012 8480 6040 8588
rect 6457 8585 6469 8588
rect 6503 8585 6515 8619
rect 6457 8579 6515 8585
rect 7098 8576 7104 8628
rect 7156 8576 7162 8628
rect 7193 8619 7251 8625
rect 7193 8585 7205 8619
rect 7239 8585 7251 8619
rect 7193 8579 7251 8585
rect 6825 8551 6883 8557
rect 6825 8517 6837 8551
rect 6871 8548 6883 8551
rect 7009 8551 7067 8557
rect 7009 8548 7021 8551
rect 6871 8520 7021 8548
rect 6871 8517 6883 8520
rect 6825 8511 6883 8517
rect 7009 8517 7021 8520
rect 7055 8517 7067 8551
rect 7009 8511 7067 8517
rect 5592 8452 6040 8480
rect 5592 8440 5598 8452
rect 6362 8440 6368 8492
rect 6420 8440 6426 8492
rect 6638 8440 6644 8492
rect 6696 8440 6702 8492
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8480 6975 8483
rect 7116 8480 7144 8576
rect 7208 8548 7236 8579
rect 7466 8576 7472 8628
rect 7524 8616 7530 8628
rect 7650 8616 7656 8628
rect 7524 8588 7656 8616
rect 7524 8576 7530 8588
rect 7650 8576 7656 8588
rect 7708 8616 7714 8628
rect 8941 8619 8999 8625
rect 8941 8616 8953 8619
rect 7708 8588 8953 8616
rect 7708 8576 7714 8588
rect 8941 8585 8953 8588
rect 8987 8585 8999 8619
rect 8941 8579 8999 8585
rect 7806 8551 7864 8557
rect 7806 8548 7818 8551
rect 7208 8520 7818 8548
rect 7806 8517 7818 8520
rect 7852 8517 7864 8551
rect 7806 8511 7864 8517
rect 6963 8452 7144 8480
rect 6963 8449 6975 8452
rect 6917 8443 6975 8449
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8480 7527 8483
rect 7650 8480 7656 8492
rect 7515 8452 7656 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 4522 8412 4528 8424
rect 3804 8384 4528 8412
rect 4522 8372 4528 8384
rect 4580 8372 4586 8424
rect 6380 8412 6408 8440
rect 6380 8384 6684 8412
rect 4246 8304 4252 8356
rect 4304 8344 4310 8356
rect 5258 8344 5264 8356
rect 4304 8316 5264 8344
rect 4304 8304 4310 8316
rect 5258 8304 5264 8316
rect 5316 8344 5322 8356
rect 6380 8344 6408 8384
rect 6656 8356 6684 8384
rect 7374 8372 7380 8424
rect 7432 8412 7438 8424
rect 7561 8415 7619 8421
rect 7561 8412 7573 8415
rect 7432 8384 7573 8412
rect 7432 8372 7438 8384
rect 7561 8381 7573 8384
rect 7607 8381 7619 8415
rect 7561 8375 7619 8381
rect 5316 8316 6408 8344
rect 5316 8304 5322 8316
rect 6638 8304 6644 8356
rect 6696 8304 6702 8356
rect 3108 8248 3372 8276
rect 3108 8236 3114 8248
rect 3878 8236 3884 8288
rect 3936 8236 3942 8288
rect 5350 8236 5356 8288
rect 5408 8276 5414 8288
rect 6270 8276 6276 8288
rect 5408 8248 6276 8276
rect 5408 8236 5414 8248
rect 6270 8236 6276 8248
rect 6328 8276 6334 8288
rect 6730 8276 6736 8288
rect 6328 8248 6736 8276
rect 6328 8236 6334 8248
rect 6730 8236 6736 8248
rect 6788 8236 6794 8288
rect 1104 8186 9292 8208
rect 1104 8134 1973 8186
rect 2025 8134 2037 8186
rect 2089 8134 2101 8186
rect 2153 8134 2165 8186
rect 2217 8134 2229 8186
rect 2281 8134 4020 8186
rect 4072 8134 4084 8186
rect 4136 8134 4148 8186
rect 4200 8134 4212 8186
rect 4264 8134 4276 8186
rect 4328 8134 6067 8186
rect 6119 8134 6131 8186
rect 6183 8134 6195 8186
rect 6247 8134 6259 8186
rect 6311 8134 6323 8186
rect 6375 8134 8114 8186
rect 8166 8134 8178 8186
rect 8230 8134 8242 8186
rect 8294 8134 8306 8186
rect 8358 8134 8370 8186
rect 8422 8134 9292 8186
rect 1104 8112 9292 8134
rect 1486 8032 1492 8084
rect 1544 8072 1550 8084
rect 1765 8075 1823 8081
rect 1765 8072 1777 8075
rect 1544 8044 1777 8072
rect 1544 8032 1550 8044
rect 1765 8041 1777 8044
rect 1811 8041 1823 8075
rect 1765 8035 1823 8041
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 3326 8072 3332 8084
rect 2832 8044 3332 8072
rect 2832 8032 2838 8044
rect 3326 8032 3332 8044
rect 3384 8032 3390 8084
rect 3605 8075 3663 8081
rect 3605 8041 3617 8075
rect 3651 8072 3663 8075
rect 3878 8072 3884 8084
rect 3651 8044 3884 8072
rect 3651 8041 3663 8044
rect 3605 8035 3663 8041
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 4338 8032 4344 8084
rect 4396 8072 4402 8084
rect 5353 8075 5411 8081
rect 5353 8072 5365 8075
rect 4396 8044 5365 8072
rect 4396 8032 4402 8044
rect 5353 8041 5365 8044
rect 5399 8041 5411 8075
rect 5353 8035 5411 8041
rect 5718 8032 5724 8084
rect 5776 8032 5782 8084
rect 7190 8032 7196 8084
rect 7248 8032 7254 8084
rect 7282 8032 7288 8084
rect 7340 8032 7346 8084
rect 7466 8032 7472 8084
rect 7524 8032 7530 8084
rect 7650 8032 7656 8084
rect 7708 8072 7714 8084
rect 7745 8075 7803 8081
rect 7745 8072 7757 8075
rect 7708 8044 7757 8072
rect 7708 8032 7714 8044
rect 7745 8041 7757 8044
rect 7791 8041 7803 8075
rect 7745 8035 7803 8041
rect 1578 7964 1584 8016
rect 1636 8004 1642 8016
rect 3789 8007 3847 8013
rect 3789 8004 3801 8007
rect 1636 7976 3801 8004
rect 1636 7964 1642 7976
rect 3789 7973 3801 7976
rect 3835 7973 3847 8007
rect 3789 7967 3847 7973
rect 5902 7964 5908 8016
rect 5960 8004 5966 8016
rect 6178 8004 6184 8016
rect 5960 7976 6184 8004
rect 5960 7964 5966 7976
rect 6178 7964 6184 7976
rect 6236 8004 6242 8016
rect 6914 8004 6920 8016
rect 6236 7976 6920 8004
rect 6236 7964 6242 7976
rect 6914 7964 6920 7976
rect 6972 7964 6978 8016
rect 8018 8004 8024 8016
rect 7116 7976 8024 8004
rect 2774 7936 2780 7948
rect 2240 7908 2780 7936
rect 1762 7828 1768 7880
rect 1820 7828 1826 7880
rect 2240 7877 2268 7908
rect 2774 7896 2780 7908
rect 2832 7896 2838 7948
rect 2866 7896 2872 7948
rect 2924 7936 2930 7948
rect 3053 7939 3111 7945
rect 3053 7936 3065 7939
rect 2924 7908 3065 7936
rect 2924 7896 2930 7908
rect 3053 7905 3065 7908
rect 3099 7936 3111 7939
rect 3418 7936 3424 7948
rect 3099 7908 3424 7936
rect 3099 7905 3111 7908
rect 3053 7899 3111 7905
rect 3418 7896 3424 7908
rect 3476 7896 3482 7948
rect 4522 7896 4528 7948
rect 4580 7936 4586 7948
rect 4709 7939 4767 7945
rect 4709 7936 4721 7939
rect 4580 7908 4721 7936
rect 4580 7896 4586 7908
rect 4709 7905 4721 7908
rect 4755 7905 4767 7939
rect 4709 7899 4767 7905
rect 5074 7896 5080 7948
rect 5132 7896 5138 7948
rect 5920 7936 5948 7964
rect 6546 7936 6552 7948
rect 5644 7908 5948 7936
rect 6104 7908 6552 7936
rect 2225 7871 2283 7877
rect 2225 7837 2237 7871
rect 2271 7837 2283 7871
rect 2225 7831 2283 7837
rect 2409 7871 2467 7877
rect 2409 7837 2421 7871
rect 2455 7837 2467 7871
rect 2409 7831 2467 7837
rect 1581 7803 1639 7809
rect 1581 7769 1593 7803
rect 1627 7800 1639 7803
rect 1780 7800 1808 7828
rect 2314 7800 2320 7812
rect 1627 7772 2320 7800
rect 1627 7769 1639 7772
rect 1581 7763 1639 7769
rect 2314 7760 2320 7772
rect 2372 7760 2378 7812
rect 2424 7800 2452 7831
rect 2682 7828 2688 7880
rect 2740 7828 2746 7880
rect 2958 7828 2964 7880
rect 3016 7868 3022 7880
rect 3329 7871 3387 7877
rect 3329 7868 3341 7871
rect 3016 7840 3341 7868
rect 3016 7828 3022 7840
rect 3329 7837 3341 7840
rect 3375 7837 3387 7871
rect 3329 7831 3387 7837
rect 3602 7828 3608 7880
rect 3660 7868 3666 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3660 7840 3985 7868
rect 3660 7828 3666 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4338 7828 4344 7880
rect 4396 7868 4402 7880
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 4396 7840 5181 7868
rect 4396 7828 4402 7840
rect 5169 7837 5181 7840
rect 5215 7868 5227 7871
rect 5350 7868 5356 7880
rect 5215 7840 5356 7868
rect 5215 7837 5227 7840
rect 5169 7831 5227 7837
rect 5350 7828 5356 7840
rect 5408 7828 5414 7880
rect 5644 7877 5672 7908
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 5810 7828 5816 7880
rect 5868 7828 5874 7880
rect 5902 7828 5908 7880
rect 5960 7868 5966 7880
rect 6104 7877 6132 7908
rect 6546 7896 6552 7908
rect 6604 7936 6610 7948
rect 6604 7908 7052 7936
rect 6604 7896 6610 7908
rect 6089 7871 6147 7877
rect 6089 7868 6101 7871
rect 5960 7840 6101 7868
rect 5960 7828 5966 7840
rect 6089 7837 6101 7840
rect 6135 7837 6147 7871
rect 6089 7831 6147 7837
rect 6273 7871 6331 7877
rect 6273 7837 6285 7871
rect 6319 7837 6331 7871
rect 6273 7831 6331 7837
rect 6641 7871 6699 7877
rect 6641 7837 6653 7871
rect 6687 7837 6699 7871
rect 6641 7831 6699 7837
rect 2498 7800 2504 7812
rect 2424 7772 2504 7800
rect 2498 7760 2504 7772
rect 2556 7760 2562 7812
rect 2593 7803 2651 7809
rect 2593 7769 2605 7803
rect 2639 7800 2651 7803
rect 2639 7772 3188 7800
rect 2639 7769 2651 7772
rect 2593 7763 2651 7769
rect 1670 7692 1676 7744
rect 1728 7732 1734 7744
rect 1781 7735 1839 7741
rect 1781 7732 1793 7735
rect 1728 7704 1793 7732
rect 1728 7692 1734 7704
rect 1781 7701 1793 7704
rect 1827 7701 1839 7735
rect 1781 7695 1839 7701
rect 1949 7735 2007 7741
rect 1949 7701 1961 7735
rect 1995 7732 2007 7735
rect 2958 7732 2964 7744
rect 1995 7704 2964 7732
rect 1995 7701 2007 7704
rect 1949 7695 2007 7701
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 3160 7732 3188 7772
rect 3234 7760 3240 7812
rect 3292 7760 3298 7812
rect 5534 7800 5540 7812
rect 3344 7772 5540 7800
rect 3344 7732 3372 7772
rect 5534 7760 5540 7772
rect 5592 7760 5598 7812
rect 5718 7760 5724 7812
rect 5776 7800 5782 7812
rect 6288 7800 6316 7831
rect 5776 7772 6316 7800
rect 6656 7800 6684 7831
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 6914 7868 6920 7880
rect 6871 7840 6920 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 6914 7828 6920 7840
rect 6972 7828 6978 7880
rect 7024 7877 7052 7908
rect 7009 7871 7067 7877
rect 7009 7837 7021 7871
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 7116 7800 7144 7976
rect 8018 7964 8024 7976
rect 8076 7964 8082 8016
rect 7208 7908 7880 7936
rect 7208 7880 7236 7908
rect 7190 7828 7196 7880
rect 7248 7828 7254 7880
rect 7469 7871 7527 7877
rect 7469 7868 7481 7871
rect 7300 7840 7481 7868
rect 6656 7772 7144 7800
rect 5776 7760 5782 7772
rect 3160 7704 3372 7732
rect 3421 7735 3479 7741
rect 3421 7701 3433 7735
rect 3467 7732 3479 7735
rect 3602 7732 3608 7744
rect 3467 7704 3608 7732
rect 3467 7701 3479 7704
rect 3421 7695 3479 7701
rect 3602 7692 3608 7704
rect 3660 7732 3666 7744
rect 5810 7732 5816 7744
rect 3660 7704 5816 7732
rect 3660 7692 3666 7704
rect 5810 7692 5816 7704
rect 5868 7732 5874 7744
rect 6270 7732 6276 7744
rect 5868 7704 6276 7732
rect 5868 7692 5874 7704
rect 6270 7692 6276 7704
rect 6328 7692 6334 7744
rect 6730 7692 6736 7744
rect 6788 7732 6794 7744
rect 7300 7732 7328 7840
rect 7469 7837 7481 7840
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 7653 7871 7711 7877
rect 7653 7837 7665 7871
rect 7699 7837 7711 7871
rect 7653 7831 7711 7837
rect 6788 7704 7328 7732
rect 7668 7732 7696 7831
rect 7742 7828 7748 7880
rect 7800 7828 7806 7880
rect 7852 7877 7880 7908
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 8036 7809 8064 7964
rect 8294 7828 8300 7880
rect 8352 7828 8358 7880
rect 8021 7803 8079 7809
rect 8021 7769 8033 7803
rect 8067 7769 8079 7803
rect 8021 7763 8079 7769
rect 7742 7732 7748 7744
rect 7668 7704 7748 7732
rect 6788 7692 6794 7704
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 7926 7692 7932 7744
rect 7984 7732 7990 7744
rect 8205 7735 8263 7741
rect 8205 7732 8217 7735
rect 7984 7704 8217 7732
rect 7984 7692 7990 7704
rect 8205 7701 8217 7704
rect 8251 7701 8263 7735
rect 8205 7695 8263 7701
rect 1104 7642 9292 7664
rect 1104 7590 2633 7642
rect 2685 7590 2697 7642
rect 2749 7590 2761 7642
rect 2813 7590 2825 7642
rect 2877 7590 2889 7642
rect 2941 7590 4680 7642
rect 4732 7590 4744 7642
rect 4796 7590 4808 7642
rect 4860 7590 4872 7642
rect 4924 7590 4936 7642
rect 4988 7590 6727 7642
rect 6779 7590 6791 7642
rect 6843 7590 6855 7642
rect 6907 7590 6919 7642
rect 6971 7590 6983 7642
rect 7035 7590 8774 7642
rect 8826 7590 8838 7642
rect 8890 7590 8902 7642
rect 8954 7590 8966 7642
rect 9018 7590 9030 7642
rect 9082 7590 9292 7642
rect 1104 7568 9292 7590
rect 1302 7488 1308 7540
rect 1360 7528 1366 7540
rect 1360 7500 2360 7528
rect 1360 7488 1366 7500
rect 1394 7352 1400 7404
rect 1452 7352 1458 7404
rect 1670 7401 1676 7404
rect 1664 7355 1676 7401
rect 1670 7352 1676 7355
rect 1728 7352 1734 7404
rect 2332 7392 2360 7500
rect 2498 7488 2504 7540
rect 2556 7528 2562 7540
rect 2556 7500 2912 7528
rect 2556 7488 2562 7500
rect 2406 7420 2412 7472
rect 2464 7460 2470 7472
rect 2884 7460 2912 7500
rect 5350 7488 5356 7540
rect 5408 7488 5414 7540
rect 5626 7488 5632 7540
rect 5684 7528 5690 7540
rect 6549 7531 6607 7537
rect 6549 7528 6561 7531
rect 5684 7500 6561 7528
rect 5684 7488 5690 7500
rect 6549 7497 6561 7500
rect 6595 7497 6607 7531
rect 6549 7491 6607 7497
rect 7009 7531 7067 7537
rect 7009 7497 7021 7531
rect 7055 7528 7067 7531
rect 7558 7528 7564 7540
rect 7055 7500 7564 7528
rect 7055 7497 7067 7500
rect 7009 7491 7067 7497
rect 7558 7488 7564 7500
rect 7616 7488 7622 7540
rect 7926 7488 7932 7540
rect 7984 7488 7990 7540
rect 8205 7531 8263 7537
rect 8205 7497 8217 7531
rect 8251 7528 8263 7531
rect 8294 7528 8300 7540
rect 8251 7500 8300 7528
rect 8251 7497 8263 7500
rect 8205 7491 8263 7497
rect 8294 7488 8300 7500
rect 8352 7488 8358 7540
rect 3786 7460 3792 7472
rect 2464 7432 2774 7460
rect 2884 7432 3792 7460
rect 2464 7420 2470 7432
rect 2746 7392 2774 7432
rect 3786 7420 3792 7432
rect 3844 7460 3850 7472
rect 6089 7463 6147 7469
rect 6089 7460 6101 7463
rect 3844 7432 4108 7460
rect 3844 7420 3850 7432
rect 3605 7395 3663 7401
rect 3605 7392 3617 7395
rect 2332 7364 2452 7392
rect 2746 7364 3617 7392
rect 2424 7324 2452 7364
rect 3605 7361 3617 7364
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 2961 7327 3019 7333
rect 2961 7324 2973 7327
rect 2424 7296 2973 7324
rect 2961 7293 2973 7296
rect 3007 7293 3019 7327
rect 2961 7287 3019 7293
rect 3145 7327 3203 7333
rect 3145 7293 3157 7327
rect 3191 7293 3203 7327
rect 3145 7287 3203 7293
rect 2406 7216 2412 7268
rect 2464 7256 2470 7268
rect 2777 7259 2835 7265
rect 2777 7256 2789 7259
rect 2464 7228 2789 7256
rect 2464 7216 2470 7228
rect 2777 7225 2789 7228
rect 2823 7256 2835 7259
rect 3160 7256 3188 7287
rect 3234 7284 3240 7336
rect 3292 7284 3298 7336
rect 3326 7284 3332 7336
rect 3384 7284 3390 7336
rect 3418 7284 3424 7336
rect 3476 7284 3482 7336
rect 4080 7324 4108 7432
rect 4264 7432 4568 7460
rect 4264 7401 4292 7432
rect 4540 7404 4568 7432
rect 4724 7432 6101 7460
rect 4724 7404 4752 7432
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7361 4399 7395
rect 4341 7355 4399 7361
rect 4356 7324 4384 7355
rect 4522 7352 4528 7404
rect 4580 7352 4586 7404
rect 4706 7352 4712 7404
rect 4764 7352 4770 7404
rect 5074 7352 5080 7404
rect 5132 7352 5138 7404
rect 5258 7352 5264 7404
rect 5316 7352 5322 7404
rect 5350 7352 5356 7404
rect 5408 7352 5414 7404
rect 5828 7401 5856 7432
rect 6089 7429 6101 7432
rect 6135 7429 6147 7463
rect 6089 7423 6147 7429
rect 6380 7432 7052 7460
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7361 5687 7395
rect 5629 7355 5687 7361
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7392 6055 7395
rect 6043 7364 6132 7392
rect 6043 7361 6055 7364
rect 5997 7355 6055 7361
rect 4080 7296 4384 7324
rect 5276 7324 5304 7352
rect 5460 7324 5488 7355
rect 5276 7296 5488 7324
rect 3510 7256 3516 7268
rect 2823 7228 3516 7256
rect 2823 7225 2835 7228
rect 2777 7219 2835 7225
rect 3510 7216 3516 7228
rect 3568 7216 3574 7268
rect 4798 7216 4804 7268
rect 4856 7256 4862 7268
rect 4985 7259 5043 7265
rect 4985 7256 4997 7259
rect 4856 7228 4997 7256
rect 4856 7216 4862 7228
rect 4985 7225 4997 7228
rect 5031 7256 5043 7259
rect 5644 7256 5672 7355
rect 5031 7228 5672 7256
rect 5736 7256 5764 7355
rect 5994 7256 6000 7268
rect 5736 7228 6000 7256
rect 5031 7225 5043 7228
rect 4985 7219 5043 7225
rect 5644 7188 5672 7228
rect 5994 7216 6000 7228
rect 6052 7216 6058 7268
rect 6104 7256 6132 7364
rect 6178 7352 6184 7404
rect 6236 7352 6242 7404
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 6380 7401 6408 7432
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 6328 7364 6377 7392
rect 6328 7352 6334 7364
rect 6365 7361 6377 7364
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 6730 7352 6736 7404
rect 6788 7352 6794 7404
rect 7024 7333 7052 7432
rect 7282 7352 7288 7404
rect 7340 7352 7346 7404
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7392 7435 7395
rect 7944 7392 7972 7488
rect 7423 7364 7972 7392
rect 7423 7361 7435 7364
rect 7377 7355 7435 7361
rect 7009 7327 7067 7333
rect 7009 7293 7021 7327
rect 7055 7293 7067 7327
rect 7009 7287 7067 7293
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7293 7159 7327
rect 7101 7287 7159 7293
rect 7116 7256 7144 7287
rect 8018 7284 8024 7336
rect 8076 7284 8082 7336
rect 8754 7284 8760 7336
rect 8812 7284 8818 7336
rect 6104 7228 6592 7256
rect 6564 7200 6592 7228
rect 6656 7228 7144 7256
rect 7193 7259 7251 7265
rect 6656 7200 6684 7228
rect 7193 7225 7205 7259
rect 7239 7256 7251 7259
rect 7650 7256 7656 7268
rect 7239 7228 7656 7256
rect 7239 7225 7251 7228
rect 7193 7219 7251 7225
rect 7650 7216 7656 7228
rect 7708 7216 7714 7268
rect 6270 7188 6276 7200
rect 5644 7160 6276 7188
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 6546 7148 6552 7200
rect 6604 7148 6610 7200
rect 6638 7148 6644 7200
rect 6696 7148 6702 7200
rect 6822 7148 6828 7200
rect 6880 7148 6886 7200
rect 7466 7148 7472 7200
rect 7524 7148 7530 7200
rect 1104 7098 9292 7120
rect 1104 7046 1973 7098
rect 2025 7046 2037 7098
rect 2089 7046 2101 7098
rect 2153 7046 2165 7098
rect 2217 7046 2229 7098
rect 2281 7046 4020 7098
rect 4072 7046 4084 7098
rect 4136 7046 4148 7098
rect 4200 7046 4212 7098
rect 4264 7046 4276 7098
rect 4328 7046 6067 7098
rect 6119 7046 6131 7098
rect 6183 7046 6195 7098
rect 6247 7046 6259 7098
rect 6311 7046 6323 7098
rect 6375 7046 8114 7098
rect 8166 7046 8178 7098
rect 8230 7046 8242 7098
rect 8294 7046 8306 7098
rect 8358 7046 8370 7098
rect 8422 7046 9292 7098
rect 1104 7024 9292 7046
rect 1670 6944 1676 6996
rect 1728 6984 1734 6996
rect 1765 6987 1823 6993
rect 1765 6984 1777 6987
rect 1728 6956 1777 6984
rect 1728 6944 1734 6956
rect 1765 6953 1777 6956
rect 1811 6953 1823 6987
rect 1765 6947 1823 6953
rect 2685 6987 2743 6993
rect 2685 6953 2697 6987
rect 2731 6984 2743 6987
rect 3050 6984 3056 6996
rect 2731 6956 3056 6984
rect 2731 6953 2743 6956
rect 2685 6947 2743 6953
rect 3050 6944 3056 6956
rect 3108 6984 3114 6996
rect 3326 6984 3332 6996
rect 3108 6956 3332 6984
rect 3108 6944 3114 6956
rect 3326 6944 3332 6956
rect 3384 6984 3390 6996
rect 4062 6984 4068 6996
rect 3384 6956 4068 6984
rect 3384 6944 3390 6956
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 5350 6984 5356 6996
rect 4448 6956 5356 6984
rect 1397 6919 1455 6925
rect 1397 6885 1409 6919
rect 1443 6916 1455 6919
rect 1443 6888 1808 6916
rect 1443 6885 1455 6888
rect 1397 6879 1455 6885
rect 1486 6808 1492 6860
rect 1544 6848 1550 6860
rect 1780 6848 1808 6888
rect 2314 6876 2320 6928
rect 2372 6916 2378 6928
rect 2869 6919 2927 6925
rect 2869 6916 2881 6919
rect 2372 6888 2881 6916
rect 2372 6876 2378 6888
rect 2869 6885 2881 6888
rect 2915 6885 2927 6919
rect 2869 6879 2927 6885
rect 1949 6851 2007 6857
rect 1949 6848 1961 6851
rect 1544 6820 1716 6848
rect 1780 6820 1961 6848
rect 1544 6808 1550 6820
rect 1578 6740 1584 6792
rect 1636 6740 1642 6792
rect 1688 6789 1716 6820
rect 1949 6817 1961 6820
rect 1995 6817 2007 6851
rect 2884 6848 2912 6879
rect 3050 6848 3056 6860
rect 2884 6820 3056 6848
rect 1949 6811 2007 6817
rect 3050 6808 3056 6820
rect 3108 6808 3114 6860
rect 3326 6808 3332 6860
rect 3384 6848 3390 6860
rect 4448 6848 4476 6956
rect 5350 6944 5356 6956
rect 5408 6944 5414 6996
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 6822 6984 6828 6996
rect 5592 6956 6828 6984
rect 5592 6944 5598 6956
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 8754 6944 8760 6996
rect 8812 6944 8818 6996
rect 5258 6916 5264 6928
rect 3384 6820 3740 6848
rect 3384 6808 3390 6820
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6749 1731 6783
rect 1673 6743 1731 6749
rect 1762 6740 1768 6792
rect 1820 6740 1826 6792
rect 2038 6740 2044 6792
rect 2096 6740 2102 6792
rect 2314 6740 2320 6792
rect 2372 6780 2378 6792
rect 3142 6780 3148 6792
rect 2372 6752 3148 6780
rect 2372 6740 2378 6752
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 3234 6740 3240 6792
rect 3292 6740 3298 6792
rect 3712 6780 3740 6820
rect 4080 6820 4476 6848
rect 4540 6888 5264 6916
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 3712 6752 3801 6780
rect 3789 6749 3801 6752
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 3881 6783 3939 6789
rect 3881 6749 3893 6783
rect 3927 6780 3939 6783
rect 3970 6780 3976 6792
rect 3927 6752 3976 6780
rect 3927 6749 3939 6752
rect 3881 6743 3939 6749
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4080 6789 4108 6820
rect 4540 6792 4568 6888
rect 5258 6876 5264 6888
rect 5316 6916 5322 6928
rect 5445 6919 5503 6925
rect 5316 6888 5396 6916
rect 5316 6876 5322 6888
rect 4706 6808 4712 6860
rect 4764 6848 4770 6860
rect 4764 6820 5111 6848
rect 4764 6808 4770 6820
rect 4065 6783 4123 6789
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 4249 6783 4307 6789
rect 4249 6780 4261 6783
rect 4212 6752 4261 6780
rect 4212 6740 4218 6752
rect 4249 6749 4261 6752
rect 4295 6780 4307 6783
rect 4295 6752 4476 6780
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 1397 6715 1455 6721
rect 1397 6681 1409 6715
rect 1443 6712 1455 6715
rect 1780 6712 1808 6740
rect 2406 6712 2412 6724
rect 1443 6684 2412 6712
rect 1443 6681 1455 6684
rect 1397 6675 1455 6681
rect 2406 6672 2412 6684
rect 2464 6672 2470 6724
rect 2593 6715 2651 6721
rect 2593 6681 2605 6715
rect 2639 6712 2651 6715
rect 4338 6712 4344 6724
rect 2639 6684 4344 6712
rect 2639 6681 2651 6684
rect 2593 6675 2651 6681
rect 4338 6672 4344 6684
rect 4396 6672 4402 6724
rect 4448 6712 4476 6752
rect 4522 6740 4528 6792
rect 4580 6740 4586 6792
rect 4798 6740 4804 6792
rect 4856 6740 4862 6792
rect 4890 6740 4896 6792
rect 4948 6740 4954 6792
rect 5083 6789 5111 6820
rect 5368 6789 5396 6888
rect 5445 6885 5457 6919
rect 5491 6916 5503 6919
rect 6730 6916 6736 6928
rect 5491 6888 6316 6916
rect 5491 6885 5503 6888
rect 5445 6879 5503 6885
rect 6288 6860 6316 6888
rect 6380 6888 6736 6916
rect 6270 6808 6276 6860
rect 6328 6808 6334 6860
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 5353 6783 5411 6789
rect 5353 6749 5365 6783
rect 5399 6749 5411 6783
rect 5353 6743 5411 6749
rect 5534 6740 5540 6792
rect 5592 6780 5598 6792
rect 5721 6783 5779 6789
rect 5721 6780 5733 6783
rect 5592 6752 5733 6780
rect 5592 6740 5598 6752
rect 5721 6749 5733 6752
rect 5767 6749 5779 6783
rect 5721 6743 5779 6749
rect 6089 6783 6147 6789
rect 6089 6749 6101 6783
rect 6135 6780 6147 6783
rect 6380 6780 6408 6888
rect 6730 6876 6736 6888
rect 6788 6876 6794 6928
rect 7374 6808 7380 6860
rect 7432 6808 7438 6860
rect 6135 6752 6408 6780
rect 6135 6749 6147 6752
rect 6089 6743 6147 6749
rect 4816 6712 4844 6740
rect 4448 6684 4844 6712
rect 4982 6672 4988 6724
rect 5040 6672 5046 6724
rect 6104 6712 6132 6743
rect 6822 6740 6828 6792
rect 6880 6740 6886 6792
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6780 7067 6783
rect 7098 6780 7104 6792
rect 7055 6752 7104 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 7098 6740 7104 6752
rect 7156 6740 7162 6792
rect 7193 6783 7251 6789
rect 7193 6749 7205 6783
rect 7239 6749 7251 6783
rect 7193 6743 7251 6749
rect 7285 6783 7343 6789
rect 7285 6749 7297 6783
rect 7331 6780 7343 6783
rect 7466 6780 7472 6792
rect 7331 6752 7472 6780
rect 7331 6749 7343 6752
rect 7285 6743 7343 6749
rect 5276 6684 6132 6712
rect 3329 6647 3387 6653
rect 3329 6613 3341 6647
rect 3375 6644 3387 6647
rect 5276 6644 5304 6684
rect 6362 6672 6368 6724
rect 6420 6672 6426 6724
rect 6549 6715 6607 6721
rect 6549 6681 6561 6715
rect 6595 6712 6607 6715
rect 6840 6712 6868 6740
rect 6595 6684 6868 6712
rect 7208 6712 7236 6743
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 7650 6789 7656 6792
rect 7644 6780 7656 6789
rect 7611 6752 7656 6780
rect 7644 6743 7656 6752
rect 7650 6740 7656 6743
rect 7708 6740 7714 6792
rect 8570 6712 8576 6724
rect 7208 6684 8576 6712
rect 6595 6681 6607 6684
rect 6549 6675 6607 6681
rect 8570 6672 8576 6684
rect 8628 6672 8634 6724
rect 3375 6616 5304 6644
rect 3375 6613 3387 6616
rect 3329 6607 3387 6613
rect 5350 6604 5356 6656
rect 5408 6644 5414 6656
rect 6733 6647 6791 6653
rect 6733 6644 6745 6647
rect 5408 6616 6745 6644
rect 5408 6604 5414 6616
rect 6733 6613 6745 6616
rect 6779 6613 6791 6647
rect 6733 6607 6791 6613
rect 6825 6647 6883 6653
rect 6825 6613 6837 6647
rect 6871 6644 6883 6647
rect 7466 6644 7472 6656
rect 6871 6616 7472 6644
rect 6871 6613 6883 6616
rect 6825 6607 6883 6613
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 1104 6554 9292 6576
rect 1104 6502 2633 6554
rect 2685 6502 2697 6554
rect 2749 6502 2761 6554
rect 2813 6502 2825 6554
rect 2877 6502 2889 6554
rect 2941 6502 4680 6554
rect 4732 6502 4744 6554
rect 4796 6502 4808 6554
rect 4860 6502 4872 6554
rect 4924 6502 4936 6554
rect 4988 6502 6727 6554
rect 6779 6502 6791 6554
rect 6843 6502 6855 6554
rect 6907 6502 6919 6554
rect 6971 6502 6983 6554
rect 7035 6502 8774 6554
rect 8826 6502 8838 6554
rect 8890 6502 8902 6554
rect 8954 6502 8966 6554
rect 9018 6502 9030 6554
rect 9082 6502 9292 6554
rect 1104 6480 9292 6502
rect 1412 6412 1992 6440
rect 1412 6381 1440 6412
rect 1964 6384 1992 6412
rect 2038 6400 2044 6452
rect 2096 6400 2102 6452
rect 2133 6443 2191 6449
rect 2133 6409 2145 6443
rect 2179 6440 2191 6443
rect 2314 6440 2320 6452
rect 2179 6412 2320 6440
rect 2179 6409 2191 6412
rect 2133 6403 2191 6409
rect 2314 6400 2320 6412
rect 2372 6400 2378 6452
rect 2593 6443 2651 6449
rect 2593 6409 2605 6443
rect 2639 6440 2651 6443
rect 2866 6440 2872 6452
rect 2639 6412 2872 6440
rect 2639 6409 2651 6412
rect 2593 6403 2651 6409
rect 2866 6400 2872 6412
rect 2924 6400 2930 6452
rect 3237 6443 3295 6449
rect 3237 6409 3249 6443
rect 3283 6440 3295 6443
rect 4154 6440 4160 6452
rect 3283 6412 4160 6440
rect 3283 6409 3295 6412
rect 3237 6403 3295 6409
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 4356 6412 5488 6440
rect 1397 6375 1455 6381
rect 1397 6341 1409 6375
rect 1443 6341 1455 6375
rect 1397 6335 1455 6341
rect 1627 6341 1685 6347
rect 1627 6338 1639 6341
rect 1612 6316 1639 6338
rect 1578 6264 1584 6316
rect 1636 6307 1639 6316
rect 1673 6307 1685 6341
rect 1946 6332 1952 6384
rect 2004 6332 2010 6384
rect 2056 6372 2084 6400
rect 3510 6372 3516 6384
rect 2056 6344 3516 6372
rect 3510 6332 3516 6344
rect 3568 6332 3574 6384
rect 3786 6332 3792 6384
rect 3844 6332 3850 6384
rect 4356 6372 4384 6412
rect 4080 6344 4384 6372
rect 1636 6301 1685 6307
rect 1636 6264 1642 6301
rect 1854 6264 1860 6316
rect 1912 6304 1918 6316
rect 2225 6307 2283 6313
rect 2225 6304 2237 6307
rect 1912 6276 2237 6304
rect 1912 6264 1918 6276
rect 2225 6273 2237 6276
rect 2271 6304 2283 6307
rect 3053 6307 3111 6313
rect 3053 6304 3065 6307
rect 2271 6276 3065 6304
rect 2271 6273 2283 6276
rect 2225 6267 2283 6273
rect 3053 6273 3065 6276
rect 3099 6273 3111 6307
rect 3053 6267 3111 6273
rect 3329 6307 3387 6313
rect 3329 6273 3341 6307
rect 3375 6273 3387 6307
rect 3804 6304 3832 6332
rect 3329 6267 3387 6273
rect 3712 6276 3832 6304
rect 1670 6196 1676 6248
rect 1728 6236 1734 6248
rect 1949 6239 2007 6245
rect 1949 6236 1961 6239
rect 1728 6208 1961 6236
rect 1728 6196 1734 6208
rect 1949 6205 1961 6208
rect 1995 6205 2007 6239
rect 1949 6199 2007 6205
rect 2590 6196 2596 6248
rect 2648 6236 2654 6248
rect 2777 6239 2835 6245
rect 2777 6236 2789 6239
rect 2648 6208 2789 6236
rect 2648 6196 2654 6208
rect 2777 6205 2789 6208
rect 2823 6205 2835 6239
rect 2777 6199 2835 6205
rect 2961 6239 3019 6245
rect 2961 6205 2973 6239
rect 3007 6205 3019 6239
rect 2961 6199 3019 6205
rect 1765 6171 1823 6177
rect 1765 6137 1777 6171
rect 1811 6168 1823 6171
rect 2976 6168 3004 6199
rect 1811 6140 3004 6168
rect 3344 6168 3372 6267
rect 3418 6196 3424 6248
rect 3476 6196 3482 6248
rect 3510 6196 3516 6248
rect 3568 6196 3574 6248
rect 3712 6245 3740 6276
rect 3878 6264 3884 6316
rect 3936 6264 3942 6316
rect 3697 6239 3755 6245
rect 3697 6205 3709 6239
rect 3743 6205 3755 6239
rect 3697 6199 3755 6205
rect 3786 6196 3792 6248
rect 3844 6196 3850 6248
rect 3970 6196 3976 6248
rect 4028 6196 4034 6248
rect 3804 6168 3832 6196
rect 4080 6168 4108 6344
rect 4430 6332 4436 6384
rect 4488 6332 4494 6384
rect 5460 6372 5488 6412
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 5721 6443 5779 6449
rect 5721 6440 5733 6443
rect 5592 6412 5733 6440
rect 5592 6400 5598 6412
rect 5721 6409 5733 6412
rect 5767 6409 5779 6443
rect 6362 6440 6368 6452
rect 5721 6403 5779 6409
rect 6104 6412 6368 6440
rect 6104 6372 6132 6412
rect 6362 6400 6368 6412
rect 6420 6400 6426 6452
rect 6638 6400 6644 6452
rect 6696 6440 6702 6452
rect 6917 6443 6975 6449
rect 6917 6440 6929 6443
rect 6696 6412 6929 6440
rect 6696 6400 6702 6412
rect 6917 6409 6929 6412
rect 6963 6409 6975 6443
rect 7190 6440 7196 6452
rect 6917 6403 6975 6409
rect 7024 6412 7196 6440
rect 5460 6344 6132 6372
rect 6178 6332 6184 6384
rect 6236 6372 6242 6384
rect 6822 6372 6828 6384
rect 6236 6344 6828 6372
rect 6236 6332 6242 6344
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6273 4215 6307
rect 4157 6267 4215 6273
rect 4172 6236 4200 6267
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 5902 6304 5908 6316
rect 5592 6276 5908 6304
rect 5592 6264 5598 6276
rect 5902 6264 5908 6276
rect 5960 6264 5966 6316
rect 6564 6313 6592 6344
rect 6822 6332 6828 6344
rect 6880 6332 6886 6384
rect 7024 6316 7052 6412
rect 7190 6400 7196 6412
rect 7248 6400 7254 6452
rect 7374 6400 7380 6452
rect 7432 6400 7438 6452
rect 7466 6400 7472 6452
rect 7524 6440 7530 6452
rect 7524 6412 7604 6440
rect 7524 6400 7530 6412
rect 7392 6372 7420 6400
rect 7576 6372 7604 6412
rect 8018 6400 8024 6452
rect 8076 6440 8082 6452
rect 8754 6440 8760 6452
rect 8076 6412 8760 6440
rect 8076 6400 8082 6412
rect 8754 6400 8760 6412
rect 8812 6440 8818 6452
rect 8849 6443 8907 6449
rect 8849 6440 8861 6443
rect 8812 6412 8861 6440
rect 8812 6400 8818 6412
rect 8849 6409 8861 6412
rect 8895 6409 8907 6443
rect 8849 6403 8907 6409
rect 7714 6375 7772 6381
rect 7714 6372 7726 6375
rect 7392 6344 7512 6372
rect 7576 6344 7726 6372
rect 6457 6307 6515 6313
rect 6457 6273 6469 6307
rect 6503 6273 6515 6307
rect 6457 6267 6515 6273
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 4430 6236 4436 6248
rect 4172 6208 4436 6236
rect 4430 6196 4436 6208
rect 4488 6196 4494 6248
rect 6472 6236 6500 6267
rect 6472 6208 6592 6236
rect 6564 6180 6592 6208
rect 3344 6140 3639 6168
rect 3804 6140 4108 6168
rect 1811 6137 1823 6140
rect 1765 6131 1823 6137
rect 1486 6060 1492 6112
rect 1544 6100 1550 6112
rect 1581 6103 1639 6109
rect 1581 6100 1593 6103
rect 1544 6072 1593 6100
rect 1544 6060 1550 6072
rect 1581 6069 1593 6072
rect 1627 6069 1639 6103
rect 1581 6063 1639 6069
rect 2314 6060 2320 6112
rect 2372 6100 2378 6112
rect 3234 6100 3240 6112
rect 2372 6072 3240 6100
rect 2372 6060 2378 6072
rect 3234 6060 3240 6072
rect 3292 6060 3298 6112
rect 3611 6100 3639 6140
rect 4338 6128 4344 6180
rect 4396 6128 4402 6180
rect 6546 6128 6552 6180
rect 6604 6128 6610 6180
rect 5350 6100 5356 6112
rect 3611 6072 5356 6100
rect 5350 6060 5356 6072
rect 5408 6060 5414 6112
rect 6454 6060 6460 6112
rect 6512 6100 6518 6112
rect 6656 6100 6684 6267
rect 6748 6168 6776 6267
rect 7006 6264 7012 6316
rect 7064 6264 7070 6316
rect 7101 6307 7159 6313
rect 7101 6273 7113 6307
rect 7147 6273 7159 6307
rect 7101 6267 7159 6273
rect 6914 6196 6920 6248
rect 6972 6236 6978 6248
rect 7116 6236 7144 6267
rect 7190 6264 7196 6316
rect 7248 6264 7254 6316
rect 7484 6313 7512 6344
rect 7714 6341 7726 6344
rect 7760 6341 7772 6375
rect 7714 6335 7772 6341
rect 7377 6307 7435 6313
rect 7377 6273 7389 6307
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6273 7527 6307
rect 8018 6304 8024 6316
rect 7469 6267 7527 6273
rect 7576 6276 8024 6304
rect 7282 6236 7288 6248
rect 6972 6208 7288 6236
rect 6972 6196 6978 6208
rect 7282 6196 7288 6208
rect 7340 6196 7346 6248
rect 7392 6236 7420 6267
rect 7576 6236 7604 6276
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 7392 6208 7604 6236
rect 7466 6168 7472 6180
rect 6748 6140 7472 6168
rect 7466 6128 7472 6140
rect 7524 6128 7530 6180
rect 6512 6072 6684 6100
rect 6512 6060 6518 6072
rect 7282 6060 7288 6112
rect 7340 6060 7346 6112
rect 7374 6060 7380 6112
rect 7432 6100 7438 6112
rect 7834 6100 7840 6112
rect 7432 6072 7840 6100
rect 7432 6060 7438 6072
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 1104 6010 9292 6032
rect 1104 5958 1973 6010
rect 2025 5958 2037 6010
rect 2089 5958 2101 6010
rect 2153 5958 2165 6010
rect 2217 5958 2229 6010
rect 2281 5958 4020 6010
rect 4072 5958 4084 6010
rect 4136 5958 4148 6010
rect 4200 5958 4212 6010
rect 4264 5958 4276 6010
rect 4328 5958 6067 6010
rect 6119 5958 6131 6010
rect 6183 5958 6195 6010
rect 6247 5958 6259 6010
rect 6311 5958 6323 6010
rect 6375 5958 8114 6010
rect 8166 5958 8178 6010
rect 8230 5958 8242 6010
rect 8294 5958 8306 6010
rect 8358 5958 8370 6010
rect 8422 5958 9292 6010
rect 1104 5936 9292 5958
rect 3142 5856 3148 5908
rect 3200 5856 3206 5908
rect 3326 5856 3332 5908
rect 3384 5896 3390 5908
rect 3510 5896 3516 5908
rect 3384 5868 3516 5896
rect 3384 5856 3390 5868
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 4338 5856 4344 5908
rect 4396 5896 4402 5908
rect 4396 5868 5028 5896
rect 4396 5856 4402 5868
rect 2777 5831 2835 5837
rect 2777 5797 2789 5831
rect 2823 5828 2835 5831
rect 3786 5828 3792 5840
rect 2823 5800 3792 5828
rect 2823 5797 2835 5800
rect 2777 5791 2835 5797
rect 3786 5788 3792 5800
rect 3844 5828 3850 5840
rect 5000 5837 5028 5868
rect 5074 5856 5080 5908
rect 5132 5896 5138 5908
rect 5169 5899 5227 5905
rect 5169 5896 5181 5899
rect 5132 5868 5181 5896
rect 5132 5856 5138 5868
rect 5169 5865 5181 5868
rect 5215 5865 5227 5899
rect 5169 5859 5227 5865
rect 5353 5899 5411 5905
rect 5353 5865 5365 5899
rect 5399 5896 5411 5899
rect 5718 5896 5724 5908
rect 5399 5868 5724 5896
rect 5399 5865 5411 5868
rect 5353 5859 5411 5865
rect 5718 5856 5724 5868
rect 5776 5856 5782 5908
rect 6457 5899 6515 5905
rect 6457 5865 6469 5899
rect 6503 5896 6515 5899
rect 7098 5896 7104 5908
rect 6503 5868 7104 5896
rect 6503 5865 6515 5868
rect 6457 5859 6515 5865
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 7466 5856 7472 5908
rect 7524 5856 7530 5908
rect 8202 5856 8208 5908
rect 8260 5856 8266 5908
rect 4985 5831 5043 5837
rect 3844 5800 4752 5828
rect 3844 5788 3850 5800
rect 2406 5720 2412 5772
rect 2464 5760 2470 5772
rect 3234 5760 3240 5772
rect 2464 5732 3240 5760
rect 2464 5720 2470 5732
rect 3234 5720 3240 5732
rect 3292 5760 3298 5772
rect 3292 5732 3464 5760
rect 3292 5720 3298 5732
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 1664 5695 1722 5701
rect 1664 5661 1676 5695
rect 1710 5692 1722 5695
rect 2590 5692 2596 5704
rect 1710 5664 2596 5692
rect 1710 5661 1722 5664
rect 1664 5655 1722 5661
rect 2590 5652 2596 5664
rect 2648 5652 2654 5704
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5692 2927 5695
rect 3329 5695 3387 5701
rect 3329 5692 3341 5695
rect 2915 5664 3341 5692
rect 2915 5661 2927 5664
rect 2869 5655 2927 5661
rect 3329 5661 3341 5664
rect 3375 5661 3387 5695
rect 3436 5692 3464 5732
rect 3510 5720 3516 5772
rect 3568 5720 3574 5772
rect 4341 5763 4399 5769
rect 3620 5732 4200 5760
rect 3620 5701 3648 5732
rect 3605 5695 3663 5701
rect 3605 5692 3617 5695
rect 3436 5664 3617 5692
rect 3329 5655 3387 5661
rect 3605 5661 3617 5664
rect 3651 5661 3663 5695
rect 3605 5655 3663 5661
rect 2498 5584 2504 5636
rect 2556 5624 2562 5636
rect 2884 5624 2912 5655
rect 2556 5596 2912 5624
rect 3344 5624 3372 5655
rect 4062 5652 4068 5704
rect 4120 5652 4126 5704
rect 4080 5624 4108 5652
rect 3344 5596 4108 5624
rect 2556 5584 2562 5596
rect 2961 5559 3019 5565
rect 2961 5525 2973 5559
rect 3007 5556 3019 5559
rect 3602 5556 3608 5568
rect 3007 5528 3608 5556
rect 3007 5525 3019 5528
rect 2961 5519 3019 5525
rect 3602 5516 3608 5528
rect 3660 5516 3666 5568
rect 4172 5556 4200 5732
rect 4341 5729 4353 5763
rect 4387 5760 4399 5763
rect 4522 5760 4528 5772
rect 4387 5732 4528 5760
rect 4387 5729 4399 5732
rect 4341 5723 4399 5729
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 4724 5769 4752 5800
rect 4985 5797 4997 5831
rect 5031 5797 5043 5831
rect 4985 5791 5043 5797
rect 5258 5788 5264 5840
rect 5316 5828 5322 5840
rect 6546 5828 6552 5840
rect 5316 5800 6552 5828
rect 5316 5788 5322 5800
rect 5644 5769 5672 5800
rect 6546 5788 6552 5800
rect 6604 5828 6610 5840
rect 8220 5828 8248 5856
rect 6604 5800 8248 5828
rect 6604 5788 6610 5800
rect 8662 5788 8668 5840
rect 8720 5788 8726 5840
rect 4709 5763 4767 5769
rect 4709 5729 4721 5763
rect 4755 5729 4767 5763
rect 4709 5723 4767 5729
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5729 5687 5763
rect 5629 5723 5687 5729
rect 5718 5720 5724 5772
rect 5776 5720 5782 5772
rect 5813 5763 5871 5769
rect 5813 5729 5825 5763
rect 5859 5760 5871 5763
rect 6730 5760 6736 5772
rect 5859 5732 6736 5760
rect 5859 5729 5871 5732
rect 5813 5723 5871 5729
rect 6288 5704 6316 5732
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 7282 5720 7288 5772
rect 7340 5720 7346 5772
rect 7466 5720 7472 5772
rect 7524 5760 7530 5772
rect 7745 5763 7803 5769
rect 7745 5760 7757 5763
rect 7524 5732 7757 5760
rect 7524 5720 7530 5732
rect 7745 5729 7757 5732
rect 7791 5729 7803 5763
rect 7745 5723 7803 5729
rect 8018 5720 8024 5772
rect 8076 5760 8082 5772
rect 8680 5760 8708 5788
rect 8076 5732 8708 5760
rect 8076 5720 8082 5732
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5692 4307 5695
rect 4617 5695 4675 5701
rect 4295 5664 4568 5692
rect 4295 5661 4307 5664
rect 4249 5655 4307 5661
rect 4540 5633 4568 5664
rect 4617 5661 4629 5695
rect 4663 5692 4675 5695
rect 5074 5692 5080 5704
rect 4663 5664 5080 5692
rect 4663 5661 4675 5664
rect 4617 5655 4675 5661
rect 5074 5652 5080 5664
rect 5132 5652 5138 5704
rect 5350 5652 5356 5704
rect 5408 5692 5414 5704
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 5408 5664 5457 5692
rect 5408 5652 5414 5664
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 5902 5692 5908 5704
rect 5445 5655 5503 5661
rect 5644 5664 5908 5692
rect 4525 5627 4583 5633
rect 4525 5593 4537 5627
rect 4571 5624 4583 5627
rect 5534 5624 5540 5636
rect 4571 5596 5540 5624
rect 4571 5593 4583 5596
rect 4525 5587 4583 5593
rect 5534 5584 5540 5596
rect 5592 5584 5598 5636
rect 5644 5556 5672 5664
rect 5902 5652 5908 5664
rect 5960 5652 5966 5704
rect 6270 5652 6276 5704
rect 6328 5652 6334 5704
rect 6362 5652 6368 5704
rect 6420 5652 6426 5704
rect 6454 5652 6460 5704
rect 6512 5652 6518 5704
rect 6546 5652 6552 5704
rect 6604 5692 6610 5704
rect 6641 5695 6699 5701
rect 6641 5692 6653 5695
rect 6604 5664 6653 5692
rect 6604 5652 6610 5664
rect 6641 5661 6653 5664
rect 6687 5692 6699 5695
rect 6822 5692 6828 5704
rect 6687 5664 6828 5692
rect 6687 5661 6699 5664
rect 6641 5655 6699 5661
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 6914 5652 6920 5704
rect 6972 5652 6978 5704
rect 7006 5652 7012 5704
rect 7064 5652 7070 5704
rect 7300 5692 7328 5720
rect 7377 5695 7435 5701
rect 7377 5692 7389 5695
rect 7300 5664 7389 5692
rect 7377 5661 7389 5664
rect 7423 5661 7435 5695
rect 7377 5655 7435 5661
rect 8110 5652 8116 5704
rect 8168 5652 8174 5704
rect 8404 5701 8432 5732
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5661 8447 5695
rect 8665 5695 8723 5701
rect 8665 5692 8677 5695
rect 8389 5655 8447 5661
rect 8496 5664 8677 5692
rect 6380 5624 6408 5652
rect 5736 5596 6408 5624
rect 6472 5624 6500 5652
rect 7024 5624 7052 5652
rect 6472 5596 7052 5624
rect 7628 5627 7686 5633
rect 5736 5568 5764 5596
rect 7628 5593 7640 5627
rect 7674 5624 7686 5627
rect 8205 5627 8263 5633
rect 8205 5624 8217 5627
rect 7674 5596 8217 5624
rect 7674 5593 7686 5596
rect 7628 5587 7686 5593
rect 8205 5593 8217 5596
rect 8251 5593 8263 5627
rect 8205 5587 8263 5593
rect 8496 5568 8524 5664
rect 8665 5661 8677 5664
rect 8711 5661 8723 5695
rect 8665 5655 8723 5661
rect 8754 5652 8760 5704
rect 8812 5652 8818 5704
rect 8573 5627 8631 5633
rect 8573 5593 8585 5627
rect 8619 5624 8631 5627
rect 8772 5624 8800 5652
rect 8619 5596 8800 5624
rect 8619 5593 8631 5596
rect 8573 5587 8631 5593
rect 4172 5528 5672 5556
rect 5718 5516 5724 5568
rect 5776 5516 5782 5568
rect 6089 5559 6147 5565
rect 6089 5525 6101 5559
rect 6135 5556 6147 5559
rect 6178 5556 6184 5568
rect 6135 5528 6184 5556
rect 6135 5525 6147 5528
rect 6089 5519 6147 5525
rect 6178 5516 6184 5528
rect 6236 5516 6242 5568
rect 7098 5516 7104 5568
rect 7156 5556 7162 5568
rect 7837 5559 7895 5565
rect 7837 5556 7849 5559
rect 7156 5528 7849 5556
rect 7156 5516 7162 5528
rect 7837 5525 7849 5528
rect 7883 5525 7895 5559
rect 7837 5519 7895 5525
rect 7926 5516 7932 5568
rect 7984 5556 7990 5568
rect 8478 5556 8484 5568
rect 7984 5528 8484 5556
rect 7984 5516 7990 5528
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 1104 5466 9292 5488
rect 1104 5414 2633 5466
rect 2685 5414 2697 5466
rect 2749 5414 2761 5466
rect 2813 5414 2825 5466
rect 2877 5414 2889 5466
rect 2941 5414 4680 5466
rect 4732 5414 4744 5466
rect 4796 5414 4808 5466
rect 4860 5414 4872 5466
rect 4924 5414 4936 5466
rect 4988 5414 6727 5466
rect 6779 5414 6791 5466
rect 6843 5414 6855 5466
rect 6907 5414 6919 5466
rect 6971 5414 6983 5466
rect 7035 5414 8774 5466
rect 8826 5414 8838 5466
rect 8890 5414 8902 5466
rect 8954 5414 8966 5466
rect 9018 5414 9030 5466
rect 9082 5414 9292 5466
rect 1104 5392 9292 5414
rect 3145 5355 3203 5361
rect 3145 5321 3157 5355
rect 3191 5352 3203 5355
rect 3418 5352 3424 5364
rect 3191 5324 3424 5352
rect 3191 5321 3203 5324
rect 3145 5315 3203 5321
rect 3418 5312 3424 5324
rect 3476 5312 3482 5364
rect 3510 5312 3516 5364
rect 3568 5352 3574 5364
rect 3568 5324 5672 5352
rect 3568 5312 3574 5324
rect 5644 5296 5672 5324
rect 7190 5312 7196 5364
rect 7248 5352 7254 5364
rect 7926 5352 7932 5364
rect 7248 5324 7932 5352
rect 7248 5312 7254 5324
rect 7926 5312 7932 5324
rect 7984 5312 7990 5364
rect 8018 5312 8024 5364
rect 8076 5312 8082 5364
rect 8110 5312 8116 5364
rect 8168 5312 8174 5364
rect 8202 5312 8208 5364
rect 8260 5312 8266 5364
rect 8570 5312 8576 5364
rect 8628 5352 8634 5364
rect 8665 5355 8723 5361
rect 8665 5352 8677 5355
rect 8628 5324 8677 5352
rect 8628 5312 8634 5324
rect 8665 5321 8677 5324
rect 8711 5321 8723 5355
rect 8665 5315 8723 5321
rect 2746 5256 3556 5284
rect 1394 5176 1400 5228
rect 1452 5176 1458 5228
rect 1664 5219 1722 5225
rect 1664 5185 1676 5219
rect 1710 5216 1722 5219
rect 2746 5216 2774 5256
rect 3528 5228 3556 5256
rect 3694 5244 3700 5296
rect 3752 5244 3758 5296
rect 5166 5284 5172 5296
rect 4632 5256 5172 5284
rect 1710 5188 2774 5216
rect 2961 5219 3019 5225
rect 1710 5185 1722 5188
rect 1664 5179 1722 5185
rect 2961 5185 2973 5219
rect 3007 5185 3019 5219
rect 2961 5179 3019 5185
rect 2976 5148 3004 5179
rect 3050 5176 3056 5228
rect 3108 5216 3114 5228
rect 3145 5219 3203 5225
rect 3145 5216 3157 5219
rect 3108 5188 3157 5216
rect 3108 5176 3114 5188
rect 3145 5185 3157 5188
rect 3191 5185 3203 5219
rect 3145 5179 3203 5185
rect 3510 5176 3516 5228
rect 3568 5176 3574 5228
rect 3605 5151 3663 5157
rect 3605 5148 3617 5151
rect 2976 5120 3617 5148
rect 3605 5117 3617 5120
rect 3651 5148 3663 5151
rect 3712 5148 3740 5244
rect 3786 5176 3792 5228
rect 3844 5216 3850 5228
rect 3881 5219 3939 5225
rect 3881 5216 3893 5219
rect 3844 5188 3893 5216
rect 3844 5176 3850 5188
rect 3881 5185 3893 5188
rect 3927 5185 3939 5219
rect 3881 5179 3939 5185
rect 4338 5176 4344 5228
rect 4396 5176 4402 5228
rect 4632 5225 4660 5256
rect 5166 5244 5172 5256
rect 5224 5244 5230 5296
rect 5626 5244 5632 5296
rect 5684 5284 5690 5296
rect 6454 5284 6460 5296
rect 5684 5256 6460 5284
rect 5684 5244 5690 5256
rect 6454 5244 6460 5256
rect 6512 5284 6518 5296
rect 6512 5256 6868 5284
rect 6512 5244 6518 5256
rect 6840 5228 6868 5256
rect 7466 5244 7472 5296
rect 7524 5284 7530 5296
rect 8128 5284 8156 5312
rect 7524 5256 8616 5284
rect 7524 5244 7530 5256
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5185 4675 5219
rect 4617 5179 4675 5185
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5185 4951 5219
rect 4893 5179 4951 5185
rect 3651 5120 3740 5148
rect 3651 5117 3663 5120
rect 3605 5111 3663 5117
rect 4062 5108 4068 5160
rect 4120 5148 4126 5160
rect 4522 5148 4528 5160
rect 4120 5120 4528 5148
rect 4120 5108 4126 5120
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 4908 5148 4936 5179
rect 4982 5176 4988 5228
rect 5040 5176 5046 5228
rect 5721 5219 5779 5225
rect 5721 5185 5733 5219
rect 5767 5185 5779 5219
rect 5721 5179 5779 5185
rect 5166 5148 5172 5160
rect 4908 5120 5172 5148
rect 5166 5108 5172 5120
rect 5224 5108 5230 5160
rect 5736 5148 5764 5179
rect 5810 5176 5816 5228
rect 5868 5216 5874 5228
rect 5905 5219 5963 5225
rect 5905 5216 5917 5219
rect 5868 5188 5917 5216
rect 5868 5176 5874 5188
rect 5905 5185 5917 5188
rect 5951 5185 5963 5219
rect 5905 5179 5963 5185
rect 6362 5176 6368 5228
rect 6420 5176 6426 5228
rect 6546 5176 6552 5228
rect 6604 5176 6610 5228
rect 6822 5176 6828 5228
rect 6880 5176 6886 5228
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 7101 5219 7159 5225
rect 7101 5216 7113 5219
rect 6972 5188 7113 5216
rect 6972 5176 6978 5188
rect 7101 5185 7113 5188
rect 7147 5216 7159 5219
rect 7190 5216 7196 5228
rect 7147 5188 7196 5216
rect 7147 5185 7159 5188
rect 7101 5179 7159 5185
rect 7190 5176 7196 5188
rect 7248 5176 7254 5228
rect 7285 5219 7343 5225
rect 7285 5185 7297 5219
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 7745 5219 7803 5225
rect 7745 5185 7757 5219
rect 7791 5216 7803 5219
rect 7834 5216 7840 5228
rect 7791 5188 7840 5216
rect 7791 5185 7803 5188
rect 7745 5179 7803 5185
rect 7006 5148 7012 5160
rect 5736 5120 7012 5148
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 3418 5040 3424 5092
rect 3476 5080 3482 5092
rect 5074 5080 5080 5092
rect 3476 5052 5080 5080
rect 3476 5040 3482 5052
rect 5074 5040 5080 5052
rect 5132 5080 5138 5092
rect 7300 5080 7328 5179
rect 7834 5176 7840 5188
rect 7892 5176 7898 5228
rect 8110 5176 8116 5228
rect 8168 5176 8174 5228
rect 8588 5225 8616 5256
rect 8205 5219 8263 5225
rect 8205 5185 8217 5219
rect 8251 5216 8263 5219
rect 8573 5219 8631 5225
rect 8251 5188 8432 5216
rect 8251 5185 8263 5188
rect 8205 5179 8263 5185
rect 8297 5151 8355 5157
rect 8297 5148 8309 5151
rect 5132 5052 7328 5080
rect 7484 5120 8309 5148
rect 5132 5040 5138 5052
rect 6564 5024 6592 5052
rect 2777 5015 2835 5021
rect 2777 4981 2789 5015
rect 2823 5012 2835 5015
rect 3602 5012 3608 5024
rect 2823 4984 3608 5012
rect 2823 4981 2835 4984
rect 2777 4975 2835 4981
rect 3602 4972 3608 4984
rect 3660 5012 3666 5024
rect 4430 5012 4436 5024
rect 3660 4984 4436 5012
rect 3660 4972 3666 4984
rect 4430 4972 4436 4984
rect 4488 4972 4494 5024
rect 4798 4972 4804 5024
rect 4856 5012 4862 5024
rect 5626 5012 5632 5024
rect 4856 4984 5632 5012
rect 4856 4972 4862 4984
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 5810 4972 5816 5024
rect 5868 5012 5874 5024
rect 6178 5012 6184 5024
rect 5868 4984 6184 5012
rect 5868 4972 5874 4984
rect 6178 4972 6184 4984
rect 6236 4972 6242 5024
rect 6454 4972 6460 5024
rect 6512 4972 6518 5024
rect 6546 4972 6552 5024
rect 6604 4972 6610 5024
rect 6730 4972 6736 5024
rect 6788 5012 6794 5024
rect 7484 5021 7512 5120
rect 8297 5117 8309 5120
rect 8343 5117 8355 5151
rect 8297 5111 8355 5117
rect 8404 5080 8432 5188
rect 8573 5185 8585 5219
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 8754 5176 8760 5228
rect 8812 5176 8818 5228
rect 8481 5151 8539 5157
rect 8481 5117 8493 5151
rect 8527 5117 8539 5151
rect 8481 5111 8539 5117
rect 7576 5052 8432 5080
rect 8496 5080 8524 5111
rect 8570 5080 8576 5092
rect 8496 5052 8576 5080
rect 7576 5024 7604 5052
rect 8570 5040 8576 5052
rect 8628 5040 8634 5092
rect 7469 5015 7527 5021
rect 7469 5012 7481 5015
rect 6788 4984 7481 5012
rect 6788 4972 6794 4984
rect 7469 4981 7481 4984
rect 7515 4981 7527 5015
rect 7469 4975 7527 4981
rect 7558 4972 7564 5024
rect 7616 4972 7622 5024
rect 7834 4972 7840 5024
rect 7892 4972 7898 5024
rect 1104 4922 9292 4944
rect 1104 4870 1973 4922
rect 2025 4870 2037 4922
rect 2089 4870 2101 4922
rect 2153 4870 2165 4922
rect 2217 4870 2229 4922
rect 2281 4870 4020 4922
rect 4072 4870 4084 4922
rect 4136 4870 4148 4922
rect 4200 4870 4212 4922
rect 4264 4870 4276 4922
rect 4328 4870 6067 4922
rect 6119 4870 6131 4922
rect 6183 4870 6195 4922
rect 6247 4870 6259 4922
rect 6311 4870 6323 4922
rect 6375 4870 8114 4922
rect 8166 4870 8178 4922
rect 8230 4870 8242 4922
rect 8294 4870 8306 4922
rect 8358 4870 8370 4922
rect 8422 4870 9292 4922
rect 1104 4848 9292 4870
rect 1578 4768 1584 4820
rect 1636 4808 1642 4820
rect 1673 4811 1731 4817
rect 1673 4808 1685 4811
rect 1636 4780 1685 4808
rect 1636 4768 1642 4780
rect 1673 4777 1685 4780
rect 1719 4777 1731 4811
rect 1673 4771 1731 4777
rect 2498 4768 2504 4820
rect 2556 4768 2562 4820
rect 2777 4811 2835 4817
rect 2777 4777 2789 4811
rect 2823 4808 2835 4811
rect 4890 4808 4896 4820
rect 2823 4780 4896 4808
rect 2823 4777 2835 4780
rect 2777 4771 2835 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 5258 4768 5264 4820
rect 5316 4808 5322 4820
rect 5718 4808 5724 4820
rect 5316 4780 5724 4808
rect 5316 4768 5322 4780
rect 5718 4768 5724 4780
rect 5776 4768 5782 4820
rect 6181 4811 6239 4817
rect 6181 4777 6193 4811
rect 6227 4808 6239 4811
rect 7466 4808 7472 4820
rect 6227 4780 7472 4808
rect 6227 4777 6239 4780
rect 6181 4771 6239 4777
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 8570 4768 8576 4820
rect 8628 4768 8634 4820
rect 2516 4740 2544 4768
rect 3418 4740 3424 4752
rect 2148 4712 2544 4740
rect 2746 4712 3424 4740
rect 1578 4564 1584 4616
rect 1636 4604 1642 4616
rect 2148 4613 2176 4712
rect 2746 4672 2774 4712
rect 3418 4700 3424 4712
rect 3476 4700 3482 4752
rect 4246 4700 4252 4752
rect 4304 4740 4310 4752
rect 5537 4743 5595 4749
rect 5537 4740 5549 4743
rect 4304 4712 5549 4740
rect 4304 4700 4310 4712
rect 5537 4709 5549 4712
rect 5583 4740 5595 4743
rect 6914 4740 6920 4752
rect 5583 4712 6920 4740
rect 5583 4709 5595 4712
rect 5537 4703 5595 4709
rect 6914 4700 6920 4712
rect 6972 4700 6978 4752
rect 8588 4740 8616 4768
rect 7024 4712 8616 4740
rect 2516 4644 2774 4672
rect 1857 4607 1915 4613
rect 1857 4604 1869 4607
rect 1636 4576 1869 4604
rect 1636 4564 1642 4576
rect 1857 4573 1869 4576
rect 1903 4604 1915 4607
rect 2133 4607 2191 4613
rect 2133 4604 2145 4607
rect 1903 4576 2145 4604
rect 1903 4573 1915 4576
rect 1857 4567 1915 4573
rect 2133 4573 2145 4576
rect 2179 4573 2191 4607
rect 2133 4567 2191 4573
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4604 2375 4607
rect 2406 4604 2412 4616
rect 2363 4576 2412 4604
rect 2363 4573 2375 4576
rect 2317 4567 2375 4573
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 2516 4613 2544 4644
rect 3142 4632 3148 4684
rect 3200 4632 3206 4684
rect 3973 4675 4031 4681
rect 3973 4672 3985 4675
rect 3712 4644 3985 4672
rect 3712 4616 3740 4644
rect 3973 4641 3985 4644
rect 4019 4641 4031 4675
rect 5077 4675 5135 4681
rect 5077 4672 5089 4675
rect 3973 4635 4031 4641
rect 4172 4644 4844 4672
rect 3602 4613 3608 4616
rect 2501 4607 2559 4613
rect 2501 4573 2513 4607
rect 2547 4573 2559 4607
rect 2501 4567 2559 4573
rect 2593 4607 2651 4613
rect 2593 4573 2605 4607
rect 2639 4573 2651 4607
rect 2593 4567 2651 4573
rect 3559 4607 3608 4613
rect 3559 4573 3571 4607
rect 3605 4573 3608 4607
rect 3559 4567 3608 4573
rect 2222 4496 2228 4548
rect 2280 4536 2286 4548
rect 2608 4536 2636 4567
rect 3602 4564 3608 4567
rect 3660 4564 3666 4616
rect 3694 4564 3700 4616
rect 3752 4564 3758 4616
rect 3786 4564 3792 4616
rect 3844 4606 3850 4616
rect 3881 4607 3939 4613
rect 3881 4606 3893 4607
rect 3844 4578 3893 4606
rect 3844 4564 3850 4578
rect 3881 4573 3893 4578
rect 3927 4573 3939 4607
rect 3881 4567 3939 4573
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4604 4123 4607
rect 4172 4604 4200 4644
rect 4816 4616 4844 4644
rect 4908 4644 5089 4672
rect 4908 4616 4936 4644
rect 5077 4641 5089 4644
rect 5123 4641 5135 4675
rect 5077 4635 5135 4641
rect 5169 4675 5227 4681
rect 5169 4641 5181 4675
rect 5215 4672 5227 4675
rect 5258 4672 5264 4684
rect 5215 4644 5264 4672
rect 5215 4641 5227 4644
rect 5169 4635 5227 4641
rect 5258 4632 5264 4644
rect 5316 4632 5322 4684
rect 5350 4632 5356 4684
rect 5408 4632 5414 4684
rect 5626 4632 5632 4684
rect 5684 4632 5690 4684
rect 7024 4672 7052 4712
rect 7834 4672 7840 4684
rect 5828 4644 7052 4672
rect 7208 4644 7840 4672
rect 4111 4576 4200 4604
rect 4249 4607 4307 4613
rect 4111 4573 4123 4576
rect 4065 4567 4123 4573
rect 4249 4573 4261 4607
rect 4295 4604 4307 4607
rect 4430 4606 4436 4616
rect 4356 4604 4436 4606
rect 4295 4578 4436 4604
rect 4295 4576 4384 4578
rect 4295 4573 4307 4576
rect 4249 4567 4307 4573
rect 4430 4564 4436 4578
rect 4488 4564 4494 4616
rect 4617 4607 4675 4613
rect 4617 4573 4629 4607
rect 4663 4573 4675 4607
rect 4617 4567 4675 4573
rect 4632 4536 4660 4567
rect 4798 4564 4804 4616
rect 4856 4564 4862 4616
rect 4890 4564 4896 4616
rect 4948 4564 4954 4616
rect 4982 4564 4988 4616
rect 5040 4564 5046 4616
rect 5184 4576 5672 4604
rect 5184 4536 5212 4576
rect 2280 4508 5212 4536
rect 5261 4539 5319 4545
rect 2280 4496 2286 4508
rect 5261 4505 5273 4539
rect 5307 4536 5319 4539
rect 5644 4536 5672 4576
rect 5718 4564 5724 4616
rect 5776 4604 5782 4616
rect 5828 4613 5856 4644
rect 5813 4607 5871 4613
rect 5813 4604 5825 4607
rect 5776 4576 5825 4604
rect 5776 4564 5782 4576
rect 5813 4573 5825 4576
rect 5859 4573 5871 4607
rect 5813 4567 5871 4573
rect 5905 4607 5963 4613
rect 5905 4573 5917 4607
rect 5951 4573 5963 4607
rect 5905 4567 5963 4573
rect 5920 4536 5948 4567
rect 5994 4564 6000 4616
rect 6052 4564 6058 4616
rect 6638 4604 6644 4616
rect 6104 4576 6644 4604
rect 6104 4536 6132 4576
rect 6638 4564 6644 4576
rect 6696 4564 6702 4616
rect 7006 4564 7012 4616
rect 7064 4604 7070 4616
rect 7208 4613 7236 4644
rect 7834 4632 7840 4644
rect 7892 4632 7898 4684
rect 7926 4632 7932 4684
rect 7984 4632 7990 4684
rect 7101 4607 7159 4613
rect 7101 4604 7113 4607
rect 7064 4576 7113 4604
rect 7064 4564 7070 4576
rect 7101 4573 7113 4576
rect 7147 4573 7159 4607
rect 7101 4567 7159 4573
rect 7193 4607 7251 4613
rect 7193 4573 7205 4607
rect 7239 4573 7251 4607
rect 7193 4567 7251 4573
rect 6457 4539 6515 4545
rect 6457 4536 6469 4539
rect 5307 4508 5396 4536
rect 5644 4508 6132 4536
rect 6196 4508 6469 4536
rect 5307 4505 5319 4508
rect 5261 4499 5319 4505
rect 1949 4471 2007 4477
rect 1949 4437 1961 4471
rect 1995 4468 2007 4471
rect 4154 4468 4160 4480
rect 1995 4440 4160 4468
rect 1995 4437 2007 4440
rect 1949 4431 2007 4437
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 4249 4471 4307 4477
rect 4249 4437 4261 4471
rect 4295 4468 4307 4471
rect 4338 4468 4344 4480
rect 4295 4440 4344 4468
rect 4295 4437 4307 4440
rect 4249 4431 4307 4437
rect 4338 4428 4344 4440
rect 4396 4428 4402 4480
rect 5368 4468 5396 4508
rect 5626 4468 5632 4480
rect 5368 4440 5632 4468
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 5994 4428 6000 4480
rect 6052 4468 6058 4480
rect 6196 4468 6224 4508
rect 6457 4505 6469 4508
rect 6503 4536 6515 4539
rect 6730 4536 6736 4548
rect 6503 4508 6736 4536
rect 6503 4505 6515 4508
rect 6457 4499 6515 4505
rect 6730 4496 6736 4508
rect 6788 4496 6794 4548
rect 7116 4536 7144 4567
rect 7282 4564 7288 4616
rect 7340 4564 7346 4616
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4604 7435 4607
rect 7466 4604 7472 4616
rect 7423 4576 7472 4604
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 7561 4607 7619 4613
rect 7561 4573 7573 4607
rect 7607 4604 7619 4607
rect 7944 4604 7972 4632
rect 7607 4576 7972 4604
rect 7607 4573 7619 4576
rect 7561 4567 7619 4573
rect 8018 4564 8024 4616
rect 8076 4564 8082 4616
rect 8205 4607 8263 4613
rect 8205 4573 8217 4607
rect 8251 4573 8263 4607
rect 8205 4567 8263 4573
rect 7837 4539 7895 4545
rect 7837 4536 7849 4539
rect 7116 4508 7849 4536
rect 7837 4505 7849 4508
rect 7883 4505 7895 4539
rect 7837 4499 7895 4505
rect 6052 4440 6224 4468
rect 6052 4428 6058 4440
rect 6270 4428 6276 4480
rect 6328 4428 6334 4480
rect 6917 4471 6975 4477
rect 6917 4437 6929 4471
rect 6963 4468 6975 4471
rect 7190 4468 7196 4480
rect 6963 4440 7196 4468
rect 6963 4437 6975 4440
rect 6917 4431 6975 4437
rect 7190 4428 7196 4440
rect 7248 4428 7254 4480
rect 7742 4428 7748 4480
rect 7800 4468 7806 4480
rect 8220 4468 8248 4567
rect 8478 4564 8484 4616
rect 8536 4564 8542 4616
rect 8294 4468 8300 4480
rect 7800 4440 8300 4468
rect 7800 4428 7806 4440
rect 8294 4428 8300 4440
rect 8352 4428 8358 4480
rect 1104 4378 9292 4400
rect 1104 4326 2633 4378
rect 2685 4326 2697 4378
rect 2749 4326 2761 4378
rect 2813 4326 2825 4378
rect 2877 4326 2889 4378
rect 2941 4326 4680 4378
rect 4732 4326 4744 4378
rect 4796 4326 4808 4378
rect 4860 4326 4872 4378
rect 4924 4326 4936 4378
rect 4988 4326 6727 4378
rect 6779 4326 6791 4378
rect 6843 4326 6855 4378
rect 6907 4326 6919 4378
rect 6971 4326 6983 4378
rect 7035 4326 8774 4378
rect 8826 4326 8838 4378
rect 8890 4326 8902 4378
rect 8954 4326 8966 4378
rect 9018 4326 9030 4378
rect 9082 4326 9292 4378
rect 1104 4304 9292 4326
rect 3694 4224 3700 4276
rect 3752 4224 3758 4276
rect 4982 4224 4988 4276
rect 5040 4264 5046 4276
rect 5258 4264 5264 4276
rect 5040 4236 5264 4264
rect 5040 4224 5046 4236
rect 5258 4224 5264 4236
rect 5316 4224 5322 4276
rect 6089 4267 6147 4273
rect 6089 4233 6101 4267
rect 6135 4264 6147 4267
rect 6454 4264 6460 4276
rect 6135 4236 6460 4264
rect 6135 4233 6147 4236
rect 6089 4227 6147 4233
rect 6454 4224 6460 4236
rect 6512 4224 6518 4276
rect 7282 4224 7288 4276
rect 7340 4264 7346 4276
rect 7929 4267 7987 4273
rect 7929 4264 7941 4267
rect 7340 4236 7941 4264
rect 7340 4224 7346 4236
rect 7929 4233 7941 4236
rect 7975 4233 7987 4267
rect 7929 4227 7987 4233
rect 3712 4196 3740 4224
rect 4890 4196 4896 4208
rect 3712 4168 4896 4196
rect 4890 4156 4896 4168
rect 4948 4196 4954 4208
rect 5350 4196 5356 4208
rect 4948 4168 5356 4196
rect 4948 4156 4954 4168
rect 5350 4156 5356 4168
rect 5408 4156 5414 4208
rect 5442 4156 5448 4208
rect 5500 4156 5506 4208
rect 6822 4156 6828 4208
rect 6880 4196 6886 4208
rect 7374 4196 7380 4208
rect 6880 4168 7380 4196
rect 6880 4156 6886 4168
rect 7374 4156 7380 4168
rect 7432 4156 7438 4208
rect 1394 4088 1400 4140
rect 1452 4088 1458 4140
rect 1670 4137 1676 4140
rect 1664 4091 1676 4137
rect 1670 4088 1676 4091
rect 1728 4088 1734 4140
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 1412 3924 1440 4088
rect 3234 4020 3240 4072
rect 3292 4060 3298 4072
rect 3421 4063 3479 4069
rect 3421 4060 3433 4063
rect 3292 4032 3433 4060
rect 3292 4020 3298 4032
rect 3421 4029 3433 4032
rect 3467 4029 3479 4063
rect 5644 4060 5672 4091
rect 5810 4088 5816 4140
rect 5868 4088 5874 4140
rect 6181 4131 6239 4137
rect 6181 4097 6193 4131
rect 6227 4128 6239 4131
rect 7006 4128 7012 4140
rect 6227 4100 7012 4128
rect 6227 4097 6239 4100
rect 6181 4091 6239 4097
rect 7006 4088 7012 4100
rect 7064 4088 7070 4140
rect 7101 4131 7159 4137
rect 7101 4097 7113 4131
rect 7147 4128 7159 4131
rect 7466 4128 7472 4140
rect 7147 4100 7472 4128
rect 7147 4097 7159 4100
rect 7101 4091 7159 4097
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 7558 4088 7564 4140
rect 7616 4088 7622 4140
rect 7926 4088 7932 4140
rect 7984 4088 7990 4140
rect 8389 4131 8447 4137
rect 8389 4128 8401 4131
rect 8036 4100 8401 4128
rect 5644 4032 6592 4060
rect 3421 4023 3479 4029
rect 4157 3995 4215 4001
rect 4157 3992 4169 3995
rect 2332 3964 4169 3992
rect 2332 3924 2360 3964
rect 4157 3961 4169 3964
rect 4203 3992 4215 3995
rect 5902 3992 5908 4004
rect 4203 3964 5908 3992
rect 4203 3961 4215 3964
rect 4157 3955 4215 3961
rect 5902 3952 5908 3964
rect 5960 3952 5966 4004
rect 6564 4001 6592 4032
rect 6638 4020 6644 4072
rect 6696 4020 6702 4072
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 7374 4060 7380 4072
rect 6871 4032 7380 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 7374 4020 7380 4032
rect 7432 4020 7438 4072
rect 7576 4060 7604 4088
rect 7484 4032 7604 4060
rect 6549 3995 6607 4001
rect 6549 3961 6561 3995
rect 6595 3961 6607 3995
rect 6656 3992 6684 4020
rect 7484 3992 7512 4032
rect 6656 3964 7512 3992
rect 7944 3992 7972 4088
rect 8036 4072 8064 4100
rect 8389 4097 8401 4100
rect 8435 4097 8447 4131
rect 8389 4091 8447 4097
rect 8478 4088 8484 4140
rect 8536 4088 8542 4140
rect 8018 4020 8024 4072
rect 8076 4020 8082 4072
rect 8113 4063 8171 4069
rect 8113 4029 8125 4063
rect 8159 4029 8171 4063
rect 8113 4023 8171 4029
rect 8205 4063 8263 4069
rect 8205 4029 8217 4063
rect 8251 4029 8263 4063
rect 8205 4023 8263 4029
rect 8128 3992 8156 4023
rect 7944 3964 8156 3992
rect 8220 3992 8248 4023
rect 8294 4020 8300 4072
rect 8352 4020 8358 4072
rect 8496 3992 8524 4088
rect 8220 3964 8524 3992
rect 6549 3955 6607 3961
rect 1412 3896 2360 3924
rect 2774 3884 2780 3936
rect 2832 3884 2838 3936
rect 2866 3884 2872 3936
rect 2924 3884 2930 3936
rect 3786 3884 3792 3936
rect 3844 3924 3850 3936
rect 5258 3924 5264 3936
rect 3844 3896 5264 3924
rect 3844 3884 3850 3896
rect 5258 3884 5264 3896
rect 5316 3884 5322 3936
rect 5810 3884 5816 3936
rect 5868 3884 5874 3936
rect 6822 3884 6828 3936
rect 6880 3884 6886 3936
rect 7098 3884 7104 3936
rect 7156 3924 7162 3936
rect 7285 3927 7343 3933
rect 7285 3924 7297 3927
rect 7156 3896 7297 3924
rect 7156 3884 7162 3896
rect 7285 3893 7297 3896
rect 7331 3893 7343 3927
rect 7484 3924 7512 3964
rect 7926 3924 7932 3936
rect 7484 3896 7932 3924
rect 7285 3887 7343 3893
rect 7926 3884 7932 3896
rect 7984 3884 7990 3936
rect 1104 3834 9292 3856
rect 1104 3782 1973 3834
rect 2025 3782 2037 3834
rect 2089 3782 2101 3834
rect 2153 3782 2165 3834
rect 2217 3782 2229 3834
rect 2281 3782 4020 3834
rect 4072 3782 4084 3834
rect 4136 3782 4148 3834
rect 4200 3782 4212 3834
rect 4264 3782 4276 3834
rect 4328 3782 6067 3834
rect 6119 3782 6131 3834
rect 6183 3782 6195 3834
rect 6247 3782 6259 3834
rect 6311 3782 6323 3834
rect 6375 3782 8114 3834
rect 8166 3782 8178 3834
rect 8230 3782 8242 3834
rect 8294 3782 8306 3834
rect 8358 3782 8370 3834
rect 8422 3782 9292 3834
rect 1104 3760 9292 3782
rect 1578 3680 1584 3732
rect 1636 3680 1642 3732
rect 1670 3680 1676 3732
rect 1728 3720 1734 3732
rect 2041 3723 2099 3729
rect 2041 3720 2053 3723
rect 1728 3692 2053 3720
rect 1728 3680 1734 3692
rect 2041 3689 2053 3692
rect 2087 3689 2099 3723
rect 2041 3683 2099 3689
rect 2133 3723 2191 3729
rect 2133 3689 2145 3723
rect 2179 3720 2191 3723
rect 2498 3720 2504 3732
rect 2179 3692 2504 3720
rect 2179 3689 2191 3692
rect 2133 3683 2191 3689
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 5074 3720 5080 3732
rect 2608 3692 5080 3720
rect 2608 3652 2636 3692
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 5258 3680 5264 3732
rect 5316 3680 5322 3732
rect 5718 3680 5724 3732
rect 5776 3720 5782 3732
rect 6365 3723 6423 3729
rect 6365 3720 6377 3723
rect 5776 3692 6377 3720
rect 5776 3680 5782 3692
rect 6365 3689 6377 3692
rect 6411 3689 6423 3723
rect 6365 3683 6423 3689
rect 7006 3680 7012 3732
rect 7064 3680 7070 3732
rect 7190 3680 7196 3732
rect 7248 3680 7254 3732
rect 7374 3680 7380 3732
rect 7432 3680 7438 3732
rect 7466 3680 7472 3732
rect 7524 3720 7530 3732
rect 8113 3723 8171 3729
rect 8113 3720 8125 3723
rect 7524 3692 8125 3720
rect 7524 3680 7530 3692
rect 8113 3689 8125 3692
rect 8159 3689 8171 3723
rect 8113 3683 8171 3689
rect 8478 3680 8484 3732
rect 8536 3680 8542 3732
rect 1964 3624 2636 3652
rect 1964 3593 1992 3624
rect 3142 3612 3148 3664
rect 3200 3652 3206 3664
rect 3973 3655 4031 3661
rect 3973 3652 3985 3655
rect 3200 3624 3985 3652
rect 3200 3612 3206 3624
rect 3973 3621 3985 3624
rect 4019 3621 4031 3655
rect 3973 3615 4031 3621
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3553 2007 3587
rect 1949 3547 2007 3553
rect 2406 3544 2412 3596
rect 2464 3544 2470 3596
rect 2774 3584 2780 3596
rect 2516 3556 2780 3584
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 1360 3488 1409 3516
rect 1360 3476 1366 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3516 2283 3519
rect 2424 3516 2452 3544
rect 2516 3525 2544 3556
rect 2774 3544 2780 3556
rect 2832 3584 2838 3596
rect 3234 3584 3240 3596
rect 2832 3556 3240 3584
rect 2832 3544 2838 3556
rect 3234 3544 3240 3556
rect 3292 3544 3298 3596
rect 3786 3544 3792 3596
rect 3844 3584 3850 3596
rect 3881 3587 3939 3593
rect 3881 3584 3893 3587
rect 3844 3556 3893 3584
rect 3844 3544 3850 3556
rect 3881 3553 3893 3556
rect 3927 3553 3939 3587
rect 3881 3547 3939 3553
rect 2271 3488 2452 3516
rect 2501 3519 2559 3525
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 2501 3485 2513 3519
rect 2547 3485 2559 3519
rect 2501 3479 2559 3485
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3516 2743 3519
rect 3142 3516 3148 3528
rect 2731 3488 3148 3516
rect 2731 3485 2743 3488
rect 2685 3479 2743 3485
rect 3142 3476 3148 3488
rect 3200 3516 3206 3528
rect 3329 3519 3387 3525
rect 3329 3516 3341 3519
rect 3200 3488 3341 3516
rect 3200 3476 3206 3488
rect 3329 3485 3341 3488
rect 3375 3485 3387 3519
rect 3329 3479 3387 3485
rect 2314 3340 2320 3392
rect 2372 3340 2378 3392
rect 2774 3340 2780 3392
rect 2832 3340 2838 3392
rect 3988 3380 4016 3615
rect 4154 3612 4160 3664
rect 4212 3612 4218 3664
rect 4430 3612 4436 3664
rect 4488 3652 4494 3664
rect 4617 3655 4675 3661
rect 4617 3652 4629 3655
rect 4488 3624 4629 3652
rect 4488 3612 4494 3624
rect 4617 3621 4629 3624
rect 4663 3621 4675 3655
rect 5276 3652 5304 3680
rect 6457 3655 6515 3661
rect 4617 3615 4675 3621
rect 4816 3624 5120 3652
rect 5276 3624 5764 3652
rect 4816 3584 4844 3624
rect 4172 3556 4844 3584
rect 4172 3525 4200 3556
rect 4890 3544 4896 3596
rect 4948 3544 4954 3596
rect 5092 3584 5120 3624
rect 5092 3556 5304 3584
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3485 4215 3519
rect 4157 3479 4215 3485
rect 4338 3476 4344 3528
rect 4396 3476 4402 3528
rect 4522 3476 4528 3528
rect 4580 3476 4586 3528
rect 4706 3476 4712 3528
rect 4764 3516 4770 3528
rect 4801 3519 4859 3525
rect 4801 3516 4813 3519
rect 4764 3488 4813 3516
rect 4764 3476 4770 3488
rect 4801 3485 4813 3488
rect 4847 3485 4859 3519
rect 4801 3479 4859 3485
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3516 5043 3519
rect 5074 3516 5080 3528
rect 5031 3488 5080 3516
rect 5031 3485 5043 3488
rect 4985 3479 5043 3485
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 5169 3519 5227 3525
rect 5169 3485 5181 3519
rect 5215 3485 5227 3519
rect 5276 3516 5304 3556
rect 5445 3519 5503 3525
rect 5445 3516 5457 3519
rect 5276 3488 5457 3516
rect 5169 3479 5227 3485
rect 5445 3485 5457 3488
rect 5491 3485 5503 3519
rect 5445 3479 5503 3485
rect 4249 3451 4307 3457
rect 4249 3417 4261 3451
rect 4295 3448 4307 3451
rect 5184 3448 5212 3479
rect 4295 3420 5212 3448
rect 4295 3417 4307 3420
rect 4249 3411 4307 3417
rect 5000 3392 5028 3420
rect 5258 3408 5264 3460
rect 5316 3408 5322 3460
rect 5460 3448 5488 3479
rect 5534 3476 5540 3528
rect 5592 3516 5598 3528
rect 5629 3519 5687 3525
rect 5629 3516 5641 3519
rect 5592 3488 5641 3516
rect 5592 3476 5598 3488
rect 5629 3485 5641 3488
rect 5675 3485 5687 3519
rect 5736 3516 5764 3624
rect 6457 3621 6469 3655
rect 6503 3652 6515 3655
rect 7098 3652 7104 3664
rect 6503 3624 7104 3652
rect 6503 3621 6515 3624
rect 6457 3615 6515 3621
rect 7098 3612 7104 3624
rect 7156 3612 7162 3664
rect 7208 3584 7236 3680
rect 7392 3652 7420 3680
rect 8297 3655 8355 3661
rect 8297 3652 8309 3655
rect 7392 3624 8309 3652
rect 8297 3621 8309 3624
rect 8343 3621 8355 3655
rect 8297 3615 8355 3621
rect 6288 3556 7236 3584
rect 7653 3587 7711 3593
rect 6288 3525 6316 3556
rect 7653 3553 7665 3587
rect 7699 3584 7711 3587
rect 7742 3584 7748 3596
rect 7699 3556 7748 3584
rect 7699 3553 7711 3556
rect 7653 3547 7711 3553
rect 7742 3544 7748 3556
rect 7800 3584 7806 3596
rect 8496 3584 8524 3680
rect 7800 3556 8524 3584
rect 7800 3544 7806 3556
rect 5905 3519 5963 3525
rect 5905 3516 5917 3519
rect 5736 3488 5917 3516
rect 5629 3479 5687 3485
rect 5905 3485 5917 3488
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 6273 3519 6331 3525
rect 6273 3485 6285 3519
rect 6319 3485 6331 3519
rect 6273 3479 6331 3485
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6512 3488 6745 3516
rect 6512 3476 6518 3488
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 6733 3479 6791 3485
rect 6825 3519 6883 3525
rect 6825 3485 6837 3519
rect 6871 3516 6883 3519
rect 7374 3516 7380 3528
rect 6871 3488 7380 3516
rect 6871 3485 6883 3488
rect 6825 3479 6883 3485
rect 7374 3476 7380 3488
rect 7432 3476 7438 3528
rect 7834 3476 7840 3528
rect 7892 3476 7898 3528
rect 7926 3476 7932 3528
rect 7984 3476 7990 3528
rect 8220 3525 8248 3556
rect 8021 3519 8079 3525
rect 8021 3485 8033 3519
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3516 8263 3519
rect 8297 3519 8355 3525
rect 8297 3516 8309 3519
rect 8251 3488 8309 3516
rect 8251 3485 8263 3488
rect 8205 3479 8263 3485
rect 8297 3485 8309 3488
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 8481 3519 8539 3525
rect 8481 3485 8493 3519
rect 8527 3485 8539 3519
rect 8481 3479 8539 3485
rect 7650 3448 7656 3460
rect 5460 3420 7656 3448
rect 7650 3408 7656 3420
rect 7708 3408 7714 3460
rect 7852 3448 7880 3476
rect 8036 3448 8064 3479
rect 8496 3448 8524 3479
rect 7852 3420 8524 3448
rect 4706 3380 4712 3392
rect 3988 3352 4712 3380
rect 4706 3340 4712 3352
rect 4764 3340 4770 3392
rect 4982 3340 4988 3392
rect 5040 3340 5046 3392
rect 5077 3383 5135 3389
rect 5077 3349 5089 3383
rect 5123 3380 5135 3383
rect 5534 3380 5540 3392
rect 5123 3352 5540 3380
rect 5123 3349 5135 3352
rect 5077 3343 5135 3349
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 7668 3380 7696 3408
rect 7837 3383 7895 3389
rect 7837 3380 7849 3383
rect 7668 3352 7849 3380
rect 7837 3349 7849 3352
rect 7883 3349 7895 3383
rect 7837 3343 7895 3349
rect 1104 3290 9292 3312
rect 1104 3238 2633 3290
rect 2685 3238 2697 3290
rect 2749 3238 2761 3290
rect 2813 3238 2825 3290
rect 2877 3238 2889 3290
rect 2941 3238 4680 3290
rect 4732 3238 4744 3290
rect 4796 3238 4808 3290
rect 4860 3238 4872 3290
rect 4924 3238 4936 3290
rect 4988 3238 6727 3290
rect 6779 3238 6791 3290
rect 6843 3238 6855 3290
rect 6907 3238 6919 3290
rect 6971 3238 6983 3290
rect 7035 3238 8774 3290
rect 8826 3238 8838 3290
rect 8890 3238 8902 3290
rect 8954 3238 8966 3290
rect 9018 3238 9030 3290
rect 9082 3238 9292 3290
rect 1104 3216 9292 3238
rect 2314 3136 2320 3188
rect 2372 3176 2378 3188
rect 4065 3179 4123 3185
rect 4065 3176 4077 3179
rect 2372 3148 4077 3176
rect 2372 3136 2378 3148
rect 4065 3145 4077 3148
rect 4111 3145 4123 3179
rect 4065 3139 4123 3145
rect 4157 3179 4215 3185
rect 4157 3145 4169 3179
rect 4203 3176 4215 3179
rect 4246 3176 4252 3188
rect 4203 3148 4252 3176
rect 4203 3145 4215 3148
rect 4157 3139 4215 3145
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 4338 3136 4344 3188
rect 4396 3176 4402 3188
rect 4433 3179 4491 3185
rect 4433 3176 4445 3179
rect 4396 3148 4445 3176
rect 4396 3136 4402 3148
rect 4433 3145 4445 3148
rect 4479 3145 4491 3179
rect 4433 3139 4491 3145
rect 5810 3136 5816 3188
rect 5868 3136 5874 3188
rect 7374 3136 7380 3188
rect 7432 3176 7438 3188
rect 7929 3179 7987 3185
rect 7929 3176 7941 3179
rect 7432 3148 7941 3176
rect 7432 3136 7438 3148
rect 7929 3145 7941 3148
rect 7975 3145 7987 3179
rect 7929 3139 7987 3145
rect 3789 3111 3847 3117
rect 3789 3077 3801 3111
rect 3835 3108 3847 3111
rect 3881 3111 3939 3117
rect 3881 3108 3893 3111
rect 3835 3080 3893 3108
rect 3835 3077 3847 3080
rect 3789 3071 3847 3077
rect 3881 3077 3893 3080
rect 3927 3108 3939 3111
rect 5074 3108 5080 3120
rect 3927 3080 5080 3108
rect 3927 3077 3939 3080
rect 3881 3071 3939 3077
rect 5074 3068 5080 3080
rect 5132 3068 5138 3120
rect 5828 3108 5856 3136
rect 6610 3111 6668 3117
rect 6610 3108 6622 3111
rect 5828 3080 6622 3108
rect 6610 3077 6622 3080
rect 6656 3077 6668 3111
rect 6610 3071 6668 3077
rect 1394 3000 1400 3052
rect 1452 3040 1458 3052
rect 1854 3049 1860 3052
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 1452 3012 1593 3040
rect 1452 3000 1458 3012
rect 1581 3009 1593 3012
rect 1627 3009 1639 3043
rect 1581 3003 1639 3009
rect 1848 3003 1860 3049
rect 1854 3000 1860 3003
rect 1912 3000 1918 3052
rect 3145 3043 3203 3049
rect 3145 3009 3157 3043
rect 3191 3009 3203 3043
rect 3145 3003 3203 3009
rect 3160 2848 3188 3003
rect 3234 3000 3240 3052
rect 3292 3000 3298 3052
rect 3605 3043 3663 3049
rect 3605 3009 3617 3043
rect 3651 3040 3663 3043
rect 3694 3040 3700 3052
rect 3651 3012 3700 3040
rect 3651 3009 3663 3012
rect 3605 3003 3663 3009
rect 3694 3000 3700 3012
rect 3752 3000 3758 3052
rect 4246 3000 4252 3052
rect 4304 3000 4310 3052
rect 4338 3000 4344 3052
rect 4396 3040 4402 3052
rect 4522 3040 4528 3052
rect 4396 3012 4528 3040
rect 4396 3000 4402 3012
rect 4522 3000 4528 3012
rect 4580 3000 4586 3052
rect 5718 3000 5724 3052
rect 5776 3049 5782 3052
rect 5776 3003 5788 3049
rect 5776 3000 5782 3003
rect 5902 3000 5908 3052
rect 5960 3040 5966 3052
rect 5997 3043 6055 3049
rect 5997 3040 6009 3043
rect 5960 3012 6009 3040
rect 5960 3000 5966 3012
rect 5997 3009 6009 3012
rect 6043 3040 6055 3043
rect 6362 3040 6368 3052
rect 6043 3012 6368 3040
rect 6043 3009 6055 3012
rect 5997 3003 6055 3009
rect 6362 3000 6368 3012
rect 6420 3000 6426 3052
rect 8018 2932 8024 2984
rect 8076 2972 8082 2984
rect 8481 2975 8539 2981
rect 8481 2972 8493 2975
rect 8076 2944 8493 2972
rect 8076 2932 8082 2944
rect 8481 2941 8493 2944
rect 8527 2941 8539 2975
rect 8481 2935 8539 2941
rect 7742 2864 7748 2916
rect 7800 2864 7806 2916
rect 2961 2839 3019 2845
rect 2961 2805 2973 2839
rect 3007 2836 3019 2839
rect 3142 2836 3148 2848
rect 3007 2808 3148 2836
rect 3007 2805 3019 2808
rect 2961 2799 3019 2805
rect 3142 2796 3148 2808
rect 3200 2796 3206 2848
rect 4614 2796 4620 2848
rect 4672 2796 4678 2848
rect 1104 2746 9292 2768
rect 1104 2694 1973 2746
rect 2025 2694 2037 2746
rect 2089 2694 2101 2746
rect 2153 2694 2165 2746
rect 2217 2694 2229 2746
rect 2281 2694 4020 2746
rect 4072 2694 4084 2746
rect 4136 2694 4148 2746
rect 4200 2694 4212 2746
rect 4264 2694 4276 2746
rect 4328 2694 6067 2746
rect 6119 2694 6131 2746
rect 6183 2694 6195 2746
rect 6247 2694 6259 2746
rect 6311 2694 6323 2746
rect 6375 2694 8114 2746
rect 8166 2694 8178 2746
rect 8230 2694 8242 2746
rect 8294 2694 8306 2746
rect 8358 2694 8370 2746
rect 8422 2694 9292 2746
rect 1104 2672 9292 2694
rect 1765 2635 1823 2641
rect 1765 2601 1777 2635
rect 1811 2632 1823 2635
rect 1854 2632 1860 2644
rect 1811 2604 1860 2632
rect 1811 2601 1823 2604
rect 1765 2595 1823 2601
rect 1854 2592 1860 2604
rect 1912 2592 1918 2644
rect 2133 2635 2191 2641
rect 2133 2601 2145 2635
rect 2179 2632 2191 2635
rect 2314 2632 2320 2644
rect 2179 2604 2320 2632
rect 2179 2601 2191 2604
rect 2133 2595 2191 2601
rect 2314 2592 2320 2604
rect 2372 2592 2378 2644
rect 2406 2592 2412 2644
rect 2464 2592 2470 2644
rect 3329 2635 3387 2641
rect 3329 2601 3341 2635
rect 3375 2632 3387 2635
rect 3510 2632 3516 2644
rect 3375 2604 3516 2632
rect 3375 2601 3387 2604
rect 3329 2595 3387 2601
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 3973 2635 4031 2641
rect 3973 2601 3985 2635
rect 4019 2632 4031 2635
rect 4338 2632 4344 2644
rect 4019 2604 4344 2632
rect 4019 2601 4031 2604
rect 3973 2595 4031 2601
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 4430 2592 4436 2644
rect 4488 2592 4494 2644
rect 5626 2592 5632 2644
rect 5684 2592 5690 2644
rect 5718 2592 5724 2644
rect 5776 2592 5782 2644
rect 6181 2635 6239 2641
rect 6181 2601 6193 2635
rect 6227 2632 6239 2635
rect 6822 2632 6828 2644
rect 6227 2604 6828 2632
rect 6227 2601 6239 2604
rect 6181 2595 6239 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 8018 2592 8024 2644
rect 8076 2592 8082 2644
rect 2685 2567 2743 2573
rect 2685 2564 2697 2567
rect 1688 2536 2697 2564
rect 1688 2496 1716 2536
rect 2685 2533 2697 2536
rect 2731 2533 2743 2567
rect 2685 2527 2743 2533
rect 3694 2524 3700 2576
rect 3752 2564 3758 2576
rect 4522 2564 4528 2576
rect 3752 2536 4528 2564
rect 3752 2524 3758 2536
rect 4522 2524 4528 2536
rect 4580 2524 4586 2576
rect 5644 2564 5672 2592
rect 5813 2567 5871 2573
rect 5813 2564 5825 2567
rect 5644 2536 5825 2564
rect 5813 2533 5825 2536
rect 5859 2533 5871 2567
rect 5813 2527 5871 2533
rect 1596 2468 1716 2496
rect 1857 2499 1915 2505
rect 1596 2437 1624 2468
rect 1857 2465 1869 2499
rect 1903 2496 1915 2499
rect 2958 2496 2964 2508
rect 1903 2468 2452 2496
rect 1903 2465 1915 2468
rect 1857 2459 1915 2465
rect 1581 2431 1639 2437
rect 1581 2397 1593 2431
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2397 1731 2431
rect 1673 2391 1731 2397
rect 1688 2360 1716 2391
rect 1762 2388 1768 2440
rect 1820 2428 1826 2440
rect 2041 2431 2099 2437
rect 2041 2428 2053 2431
rect 1820 2400 2053 2428
rect 1820 2388 1826 2400
rect 2041 2397 2053 2400
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 2424 2360 2452 2468
rect 2516 2468 2964 2496
rect 2516 2437 2544 2468
rect 2958 2456 2964 2468
rect 3016 2456 3022 2508
rect 3145 2499 3203 2505
rect 3145 2465 3157 2499
rect 3191 2496 3203 2499
rect 3878 2496 3884 2508
rect 3191 2468 3884 2496
rect 3191 2465 3203 2468
rect 3145 2459 3203 2465
rect 3878 2456 3884 2468
rect 3936 2496 3942 2508
rect 4065 2499 4123 2505
rect 4065 2496 4077 2499
rect 3936 2468 4077 2496
rect 3936 2456 3942 2468
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 2774 2388 2780 2440
rect 2832 2388 2838 2440
rect 3050 2388 3056 2440
rect 3108 2388 3114 2440
rect 3234 2388 3240 2440
rect 3292 2388 3298 2440
rect 3510 2388 3516 2440
rect 3568 2388 3574 2440
rect 3694 2388 3700 2440
rect 3752 2428 3758 2440
rect 3988 2437 4016 2468
rect 4065 2465 4077 2468
rect 4111 2465 4123 2499
rect 4065 2459 4123 2465
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 3752 2400 3801 2428
rect 3752 2388 3758 2400
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2428 4307 2431
rect 4540 2428 4568 2524
rect 6638 2456 6644 2508
rect 6696 2456 6702 2508
rect 4709 2431 4767 2437
rect 4709 2428 4721 2431
rect 4295 2400 4721 2428
rect 4295 2397 4307 2400
rect 4249 2391 4307 2397
rect 4709 2397 4721 2400
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 5261 2431 5319 2437
rect 5261 2397 5273 2431
rect 5307 2428 5319 2431
rect 5353 2431 5411 2437
rect 5353 2428 5365 2431
rect 5307 2400 5365 2428
rect 5307 2397 5319 2400
rect 5261 2391 5319 2397
rect 5353 2397 5365 2400
rect 5399 2397 5411 2431
rect 5353 2391 5411 2397
rect 5442 2388 5448 2440
rect 5500 2388 5506 2440
rect 5534 2388 5540 2440
rect 5592 2428 5598 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5592 2400 5917 2428
rect 5592 2388 5598 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2397 6055 2431
rect 5997 2391 6055 2397
rect 6908 2431 6966 2437
rect 6908 2397 6920 2431
rect 6954 2428 6966 2431
rect 7190 2428 7196 2440
rect 6954 2400 7196 2428
rect 6954 2397 6966 2400
rect 6908 2391 6966 2397
rect 1688 2332 1808 2360
rect 2424 2332 2774 2360
rect 1780 2292 1808 2332
rect 2498 2292 2504 2304
rect 1780 2264 2504 2292
rect 2498 2252 2504 2264
rect 2556 2252 2562 2304
rect 2746 2292 2774 2332
rect 5166 2320 5172 2372
rect 5224 2360 5230 2372
rect 6012 2360 6040 2391
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 5224 2332 6040 2360
rect 5224 2320 5230 2332
rect 3786 2292 3792 2304
rect 2746 2264 3792 2292
rect 3786 2252 3792 2264
rect 3844 2252 3850 2304
rect 1104 2202 9292 2224
rect 1104 2150 2633 2202
rect 2685 2150 2697 2202
rect 2749 2150 2761 2202
rect 2813 2150 2825 2202
rect 2877 2150 2889 2202
rect 2941 2150 4680 2202
rect 4732 2150 4744 2202
rect 4796 2150 4808 2202
rect 4860 2150 4872 2202
rect 4924 2150 4936 2202
rect 4988 2150 6727 2202
rect 6779 2150 6791 2202
rect 6843 2150 6855 2202
rect 6907 2150 6919 2202
rect 6971 2150 6983 2202
rect 7035 2150 8774 2202
rect 8826 2150 8838 2202
rect 8890 2150 8902 2202
rect 8954 2150 8966 2202
rect 9018 2150 9030 2202
rect 9082 2150 9292 2202
rect 1104 2128 9292 2150
<< via1 >>
rect 1973 10310 2025 10362
rect 2037 10310 2089 10362
rect 2101 10310 2153 10362
rect 2165 10310 2217 10362
rect 2229 10310 2281 10362
rect 4020 10310 4072 10362
rect 4084 10310 4136 10362
rect 4148 10310 4200 10362
rect 4212 10310 4264 10362
rect 4276 10310 4328 10362
rect 6067 10310 6119 10362
rect 6131 10310 6183 10362
rect 6195 10310 6247 10362
rect 6259 10310 6311 10362
rect 6323 10310 6375 10362
rect 8114 10310 8166 10362
rect 8178 10310 8230 10362
rect 8242 10310 8294 10362
rect 8306 10310 8358 10362
rect 8370 10310 8422 10362
rect 5816 10208 5868 10260
rect 5356 10140 5408 10192
rect 7656 10183 7708 10192
rect 7656 10149 7665 10183
rect 7665 10149 7699 10183
rect 7699 10149 7708 10183
rect 7656 10140 7708 10149
rect 7288 10072 7340 10124
rect 2044 10004 2096 10056
rect 2964 10004 3016 10056
rect 3240 10004 3292 10056
rect 5264 10004 5316 10056
rect 7196 10004 7248 10056
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 6184 9936 6236 9988
rect 7104 9936 7156 9988
rect 7472 9979 7524 9988
rect 7472 9945 7481 9979
rect 7481 9945 7515 9979
rect 7515 9945 7524 9979
rect 7472 9936 7524 9945
rect 2504 9911 2556 9920
rect 2504 9877 2513 9911
rect 2513 9877 2547 9911
rect 2547 9877 2556 9911
rect 2504 9868 2556 9877
rect 3424 9868 3476 9920
rect 4528 9868 4580 9920
rect 5080 9868 5132 9920
rect 8024 9936 8076 9988
rect 7840 9911 7892 9920
rect 7840 9877 7849 9911
rect 7849 9877 7883 9911
rect 7883 9877 7892 9911
rect 7840 9868 7892 9877
rect 2633 9766 2685 9818
rect 2697 9766 2749 9818
rect 2761 9766 2813 9818
rect 2825 9766 2877 9818
rect 2889 9766 2941 9818
rect 4680 9766 4732 9818
rect 4744 9766 4796 9818
rect 4808 9766 4860 9818
rect 4872 9766 4924 9818
rect 4936 9766 4988 9818
rect 6727 9766 6779 9818
rect 6791 9766 6843 9818
rect 6855 9766 6907 9818
rect 6919 9766 6971 9818
rect 6983 9766 7035 9818
rect 8774 9766 8826 9818
rect 8838 9766 8890 9818
rect 8902 9766 8954 9818
rect 8966 9766 9018 9818
rect 9030 9766 9082 9818
rect 1584 9707 1636 9716
rect 1584 9673 1593 9707
rect 1593 9673 1627 9707
rect 1627 9673 1636 9707
rect 1584 9664 1636 9673
rect 2044 9664 2096 9716
rect 6184 9707 6236 9716
rect 6184 9673 6193 9707
rect 6193 9673 6227 9707
rect 6227 9673 6236 9707
rect 6184 9664 6236 9673
rect 1676 9596 1728 9648
rect 1584 9528 1636 9580
rect 1584 9324 1636 9376
rect 1768 9503 1820 9512
rect 1768 9469 1777 9503
rect 1777 9469 1811 9503
rect 1811 9469 1820 9503
rect 1768 9460 1820 9469
rect 2872 9528 2924 9580
rect 4344 9528 4396 9580
rect 5724 9596 5776 9648
rect 7656 9639 7708 9648
rect 7656 9605 7690 9639
rect 7690 9605 7708 9639
rect 7656 9596 7708 9605
rect 5448 9528 5500 9580
rect 6184 9528 6236 9580
rect 7196 9571 7248 9580
rect 7196 9537 7205 9571
rect 7205 9537 7239 9571
rect 7239 9537 7248 9571
rect 7196 9528 7248 9537
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 2964 9324 3016 9376
rect 3240 9367 3292 9376
rect 3240 9333 3249 9367
rect 3249 9333 3283 9367
rect 3283 9333 3292 9367
rect 3240 9324 3292 9333
rect 4528 9324 4580 9376
rect 5540 9324 5592 9376
rect 8024 9324 8076 9376
rect 1973 9222 2025 9274
rect 2037 9222 2089 9274
rect 2101 9222 2153 9274
rect 2165 9222 2217 9274
rect 2229 9222 2281 9274
rect 4020 9222 4072 9274
rect 4084 9222 4136 9274
rect 4148 9222 4200 9274
rect 4212 9222 4264 9274
rect 4276 9222 4328 9274
rect 6067 9222 6119 9274
rect 6131 9222 6183 9274
rect 6195 9222 6247 9274
rect 6259 9222 6311 9274
rect 6323 9222 6375 9274
rect 8114 9222 8166 9274
rect 8178 9222 8230 9274
rect 8242 9222 8294 9274
rect 8306 9222 8358 9274
rect 8370 9222 8422 9274
rect 2872 9163 2924 9172
rect 2872 9129 2881 9163
rect 2881 9129 2915 9163
rect 2915 9129 2924 9163
rect 2872 9120 2924 9129
rect 5448 9120 5500 9172
rect 6000 9120 6052 9172
rect 6920 9120 6972 9172
rect 7288 9163 7340 9172
rect 7288 9129 7297 9163
rect 7297 9129 7331 9163
rect 7331 9129 7340 9163
rect 7288 9120 7340 9129
rect 7472 9120 7524 9172
rect 3148 9052 3200 9104
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 3148 8959 3200 8968
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 1492 8848 1544 8900
rect 3424 8848 3476 8900
rect 2964 8780 3016 8832
rect 3148 8780 3200 8832
rect 3884 8916 3936 8968
rect 3608 8848 3660 8900
rect 3792 8823 3844 8832
rect 3792 8789 3801 8823
rect 3801 8789 3835 8823
rect 3835 8789 3844 8823
rect 3792 8780 3844 8789
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 4252 8959 4304 8968
rect 4252 8925 4261 8959
rect 4261 8925 4295 8959
rect 4295 8925 4304 8959
rect 4252 8916 4304 8925
rect 5080 8984 5132 9036
rect 5172 8959 5224 8968
rect 5172 8925 5181 8959
rect 5181 8925 5215 8959
rect 5215 8925 5224 8959
rect 5172 8916 5224 8925
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 4620 8780 4672 8832
rect 5356 8891 5408 8900
rect 5356 8857 5387 8891
rect 5387 8857 5408 8891
rect 5356 8848 5408 8857
rect 5540 8848 5592 8900
rect 6184 8916 6236 8968
rect 6276 8916 6328 8968
rect 6644 8916 6696 8968
rect 6828 8959 6880 8968
rect 6828 8925 6837 8959
rect 6837 8925 6871 8959
rect 6871 8925 6880 8959
rect 6828 8916 6880 8925
rect 7840 8984 7892 9036
rect 7656 8959 7708 8968
rect 7656 8925 7665 8959
rect 7665 8925 7699 8959
rect 7699 8925 7708 8959
rect 7656 8916 7708 8925
rect 5816 8823 5868 8832
rect 5816 8789 5825 8823
rect 5825 8789 5859 8823
rect 5859 8789 5868 8823
rect 5816 8780 5868 8789
rect 5908 8823 5960 8832
rect 5908 8789 5917 8823
rect 5917 8789 5951 8823
rect 5951 8789 5960 8823
rect 5908 8780 5960 8789
rect 7104 8780 7156 8832
rect 7840 8780 7892 8832
rect 2633 8678 2685 8730
rect 2697 8678 2749 8730
rect 2761 8678 2813 8730
rect 2825 8678 2877 8730
rect 2889 8678 2941 8730
rect 4680 8678 4732 8730
rect 4744 8678 4796 8730
rect 4808 8678 4860 8730
rect 4872 8678 4924 8730
rect 4936 8678 4988 8730
rect 6727 8678 6779 8730
rect 6791 8678 6843 8730
rect 6855 8678 6907 8730
rect 6919 8678 6971 8730
rect 6983 8678 7035 8730
rect 8774 8678 8826 8730
rect 8838 8678 8890 8730
rect 8902 8678 8954 8730
rect 8966 8678 9018 8730
rect 9030 8678 9082 8730
rect 1492 8576 1544 8628
rect 1584 8576 1636 8628
rect 3056 8576 3108 8628
rect 1308 8440 1360 8492
rect 3148 8508 3200 8560
rect 3792 8576 3844 8628
rect 4344 8619 4396 8628
rect 4344 8585 4353 8619
rect 4353 8585 4387 8619
rect 4387 8585 4396 8619
rect 4344 8576 4396 8585
rect 5172 8576 5224 8628
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 2872 8372 2924 8424
rect 1860 8304 1912 8356
rect 3332 8440 3384 8492
rect 5908 8508 5960 8560
rect 3240 8304 3292 8356
rect 1492 8236 1544 8288
rect 1952 8236 2004 8288
rect 2964 8236 3016 8288
rect 3056 8236 3108 8288
rect 3424 8415 3476 8424
rect 3424 8381 3433 8415
rect 3433 8381 3467 8415
rect 3467 8381 3476 8415
rect 3424 8372 3476 8381
rect 3516 8415 3568 8424
rect 3516 8381 3525 8415
rect 3525 8381 3559 8415
rect 3559 8381 3568 8415
rect 3516 8372 3568 8381
rect 4344 8440 4396 8492
rect 5448 8440 5500 8492
rect 5540 8440 5592 8492
rect 7104 8576 7156 8628
rect 6368 8483 6420 8492
rect 6368 8449 6377 8483
rect 6377 8449 6411 8483
rect 6411 8449 6420 8483
rect 6368 8440 6420 8449
rect 6644 8483 6696 8492
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 7472 8576 7524 8628
rect 7656 8576 7708 8628
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 7656 8440 7708 8492
rect 4528 8372 4580 8424
rect 4252 8304 4304 8356
rect 5264 8304 5316 8356
rect 7380 8372 7432 8424
rect 6644 8304 6696 8356
rect 3884 8279 3936 8288
rect 3884 8245 3893 8279
rect 3893 8245 3927 8279
rect 3927 8245 3936 8279
rect 3884 8236 3936 8245
rect 5356 8236 5408 8288
rect 6276 8236 6328 8288
rect 6736 8236 6788 8288
rect 1973 8134 2025 8186
rect 2037 8134 2089 8186
rect 2101 8134 2153 8186
rect 2165 8134 2217 8186
rect 2229 8134 2281 8186
rect 4020 8134 4072 8186
rect 4084 8134 4136 8186
rect 4148 8134 4200 8186
rect 4212 8134 4264 8186
rect 4276 8134 4328 8186
rect 6067 8134 6119 8186
rect 6131 8134 6183 8186
rect 6195 8134 6247 8186
rect 6259 8134 6311 8186
rect 6323 8134 6375 8186
rect 8114 8134 8166 8186
rect 8178 8134 8230 8186
rect 8242 8134 8294 8186
rect 8306 8134 8358 8186
rect 8370 8134 8422 8186
rect 1492 8032 1544 8084
rect 2780 8032 2832 8084
rect 3332 8032 3384 8084
rect 3884 8032 3936 8084
rect 4344 8032 4396 8084
rect 5724 8075 5776 8084
rect 5724 8041 5733 8075
rect 5733 8041 5767 8075
rect 5767 8041 5776 8075
rect 5724 8032 5776 8041
rect 7196 8075 7248 8084
rect 7196 8041 7205 8075
rect 7205 8041 7239 8075
rect 7239 8041 7248 8075
rect 7196 8032 7248 8041
rect 7288 8075 7340 8084
rect 7288 8041 7297 8075
rect 7297 8041 7331 8075
rect 7331 8041 7340 8075
rect 7288 8032 7340 8041
rect 7472 8075 7524 8084
rect 7472 8041 7481 8075
rect 7481 8041 7515 8075
rect 7515 8041 7524 8075
rect 7472 8032 7524 8041
rect 7656 8032 7708 8084
rect 1584 7964 1636 8016
rect 5908 7964 5960 8016
rect 6184 7964 6236 8016
rect 6920 7964 6972 8016
rect 1768 7828 1820 7880
rect 2780 7896 2832 7948
rect 2872 7896 2924 7948
rect 3424 7896 3476 7948
rect 4528 7896 4580 7948
rect 5080 7939 5132 7948
rect 5080 7905 5089 7939
rect 5089 7905 5123 7939
rect 5123 7905 5132 7939
rect 5080 7896 5132 7905
rect 2320 7760 2372 7812
rect 2688 7871 2740 7880
rect 2688 7837 2697 7871
rect 2697 7837 2731 7871
rect 2731 7837 2740 7871
rect 2688 7828 2740 7837
rect 2964 7828 3016 7880
rect 3608 7828 3660 7880
rect 4344 7828 4396 7880
rect 5356 7828 5408 7880
rect 5816 7871 5868 7880
rect 5816 7837 5825 7871
rect 5825 7837 5859 7871
rect 5859 7837 5868 7871
rect 5816 7828 5868 7837
rect 5908 7828 5960 7880
rect 6552 7896 6604 7948
rect 2504 7760 2556 7812
rect 1676 7692 1728 7744
rect 2964 7692 3016 7744
rect 3240 7803 3292 7812
rect 3240 7769 3249 7803
rect 3249 7769 3283 7803
rect 3283 7769 3292 7803
rect 3240 7760 3292 7769
rect 5540 7760 5592 7812
rect 5724 7760 5776 7812
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 6920 7828 6972 7880
rect 8024 7964 8076 8016
rect 7196 7828 7248 7880
rect 3608 7692 3660 7744
rect 5816 7692 5868 7744
rect 6276 7692 6328 7744
rect 6736 7692 6788 7744
rect 7748 7871 7800 7880
rect 7748 7837 7757 7871
rect 7757 7837 7791 7871
rect 7791 7837 7800 7871
rect 7748 7828 7800 7837
rect 8300 7871 8352 7880
rect 8300 7837 8309 7871
rect 8309 7837 8343 7871
rect 8343 7837 8352 7871
rect 8300 7828 8352 7837
rect 7748 7692 7800 7744
rect 7932 7692 7984 7744
rect 2633 7590 2685 7642
rect 2697 7590 2749 7642
rect 2761 7590 2813 7642
rect 2825 7590 2877 7642
rect 2889 7590 2941 7642
rect 4680 7590 4732 7642
rect 4744 7590 4796 7642
rect 4808 7590 4860 7642
rect 4872 7590 4924 7642
rect 4936 7590 4988 7642
rect 6727 7590 6779 7642
rect 6791 7590 6843 7642
rect 6855 7590 6907 7642
rect 6919 7590 6971 7642
rect 6983 7590 7035 7642
rect 8774 7590 8826 7642
rect 8838 7590 8890 7642
rect 8902 7590 8954 7642
rect 8966 7590 9018 7642
rect 9030 7590 9082 7642
rect 1308 7488 1360 7540
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 1676 7395 1728 7404
rect 1676 7361 1710 7395
rect 1710 7361 1728 7395
rect 1676 7352 1728 7361
rect 2504 7488 2556 7540
rect 2412 7420 2464 7472
rect 5356 7531 5408 7540
rect 5356 7497 5365 7531
rect 5365 7497 5399 7531
rect 5399 7497 5408 7531
rect 5356 7488 5408 7497
rect 5632 7488 5684 7540
rect 7564 7488 7616 7540
rect 7932 7488 7984 7540
rect 8300 7488 8352 7540
rect 3792 7420 3844 7472
rect 2412 7216 2464 7268
rect 3240 7327 3292 7336
rect 3240 7293 3249 7327
rect 3249 7293 3283 7327
rect 3283 7293 3292 7327
rect 3240 7284 3292 7293
rect 3332 7327 3384 7336
rect 3332 7293 3341 7327
rect 3341 7293 3375 7327
rect 3375 7293 3384 7327
rect 3332 7284 3384 7293
rect 3424 7327 3476 7336
rect 3424 7293 3433 7327
rect 3433 7293 3467 7327
rect 3467 7293 3476 7327
rect 3424 7284 3476 7293
rect 4528 7352 4580 7404
rect 4712 7352 4764 7404
rect 5080 7395 5132 7404
rect 5080 7361 5089 7395
rect 5089 7361 5123 7395
rect 5123 7361 5132 7395
rect 5080 7352 5132 7361
rect 5264 7352 5316 7404
rect 5356 7395 5408 7404
rect 5356 7361 5365 7395
rect 5365 7361 5399 7395
rect 5399 7361 5408 7395
rect 5356 7352 5408 7361
rect 3516 7216 3568 7268
rect 4804 7216 4856 7268
rect 6000 7216 6052 7268
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 6276 7352 6328 7404
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 8024 7327 8076 7336
rect 8024 7293 8033 7327
rect 8033 7293 8067 7327
rect 8067 7293 8076 7327
rect 8024 7284 8076 7293
rect 8760 7327 8812 7336
rect 8760 7293 8769 7327
rect 8769 7293 8803 7327
rect 8803 7293 8812 7327
rect 8760 7284 8812 7293
rect 7656 7216 7708 7268
rect 6276 7148 6328 7200
rect 6552 7148 6604 7200
rect 6644 7148 6696 7200
rect 6828 7191 6880 7200
rect 6828 7157 6837 7191
rect 6837 7157 6871 7191
rect 6871 7157 6880 7191
rect 6828 7148 6880 7157
rect 7472 7191 7524 7200
rect 7472 7157 7481 7191
rect 7481 7157 7515 7191
rect 7515 7157 7524 7191
rect 7472 7148 7524 7157
rect 1973 7046 2025 7098
rect 2037 7046 2089 7098
rect 2101 7046 2153 7098
rect 2165 7046 2217 7098
rect 2229 7046 2281 7098
rect 4020 7046 4072 7098
rect 4084 7046 4136 7098
rect 4148 7046 4200 7098
rect 4212 7046 4264 7098
rect 4276 7046 4328 7098
rect 6067 7046 6119 7098
rect 6131 7046 6183 7098
rect 6195 7046 6247 7098
rect 6259 7046 6311 7098
rect 6323 7046 6375 7098
rect 8114 7046 8166 7098
rect 8178 7046 8230 7098
rect 8242 7046 8294 7098
rect 8306 7046 8358 7098
rect 8370 7046 8422 7098
rect 1676 6944 1728 6996
rect 3056 6944 3108 6996
rect 3332 6944 3384 6996
rect 4068 6944 4120 6996
rect 1492 6808 1544 6860
rect 2320 6876 2372 6928
rect 1584 6783 1636 6792
rect 1584 6749 1593 6783
rect 1593 6749 1627 6783
rect 1627 6749 1636 6783
rect 1584 6740 1636 6749
rect 3056 6808 3108 6860
rect 3332 6808 3384 6860
rect 5356 6944 5408 6996
rect 5540 6944 5592 6996
rect 6828 6944 6880 6996
rect 8760 6987 8812 6996
rect 8760 6953 8769 6987
rect 8769 6953 8803 6987
rect 8803 6953 8812 6987
rect 8760 6944 8812 6953
rect 1768 6740 1820 6792
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 2320 6783 2372 6792
rect 2320 6749 2329 6783
rect 2329 6749 2363 6783
rect 2363 6749 2372 6783
rect 2320 6740 2372 6749
rect 3148 6740 3200 6792
rect 3240 6783 3292 6792
rect 3240 6749 3249 6783
rect 3249 6749 3283 6783
rect 3283 6749 3292 6783
rect 3240 6740 3292 6749
rect 3976 6740 4028 6792
rect 5264 6876 5316 6928
rect 4712 6808 4764 6860
rect 4160 6740 4212 6792
rect 2412 6715 2464 6724
rect 2412 6681 2421 6715
rect 2421 6681 2455 6715
rect 2455 6681 2464 6715
rect 2412 6672 2464 6681
rect 4344 6672 4396 6724
rect 4528 6783 4580 6792
rect 4528 6749 4537 6783
rect 4537 6749 4571 6783
rect 4571 6749 4580 6783
rect 4528 6740 4580 6749
rect 4804 6740 4856 6792
rect 4896 6783 4948 6792
rect 4896 6749 4905 6783
rect 4905 6749 4939 6783
rect 4939 6749 4948 6783
rect 4896 6740 4948 6749
rect 6276 6808 6328 6860
rect 5540 6740 5592 6792
rect 6736 6876 6788 6928
rect 7380 6851 7432 6860
rect 7380 6817 7389 6851
rect 7389 6817 7423 6851
rect 7423 6817 7432 6851
rect 7380 6808 7432 6817
rect 4988 6715 5040 6724
rect 4988 6681 4997 6715
rect 4997 6681 5031 6715
rect 5031 6681 5040 6715
rect 4988 6672 5040 6681
rect 6828 6740 6880 6792
rect 7104 6740 7156 6792
rect 6368 6715 6420 6724
rect 6368 6681 6377 6715
rect 6377 6681 6411 6715
rect 6411 6681 6420 6715
rect 6368 6672 6420 6681
rect 7472 6740 7524 6792
rect 7656 6783 7708 6792
rect 7656 6749 7690 6783
rect 7690 6749 7708 6783
rect 7656 6740 7708 6749
rect 8576 6672 8628 6724
rect 5356 6604 5408 6656
rect 7472 6604 7524 6656
rect 2633 6502 2685 6554
rect 2697 6502 2749 6554
rect 2761 6502 2813 6554
rect 2825 6502 2877 6554
rect 2889 6502 2941 6554
rect 4680 6502 4732 6554
rect 4744 6502 4796 6554
rect 4808 6502 4860 6554
rect 4872 6502 4924 6554
rect 4936 6502 4988 6554
rect 6727 6502 6779 6554
rect 6791 6502 6843 6554
rect 6855 6502 6907 6554
rect 6919 6502 6971 6554
rect 6983 6502 7035 6554
rect 8774 6502 8826 6554
rect 8838 6502 8890 6554
rect 8902 6502 8954 6554
rect 8966 6502 9018 6554
rect 9030 6502 9082 6554
rect 2044 6400 2096 6452
rect 2320 6400 2372 6452
rect 2872 6400 2924 6452
rect 4160 6400 4212 6452
rect 1584 6264 1636 6316
rect 1952 6332 2004 6384
rect 3516 6332 3568 6384
rect 3792 6332 3844 6384
rect 1860 6264 1912 6316
rect 1676 6196 1728 6248
rect 2596 6196 2648 6248
rect 3424 6239 3476 6248
rect 3424 6205 3433 6239
rect 3433 6205 3467 6239
rect 3467 6205 3476 6239
rect 3424 6196 3476 6205
rect 3516 6239 3568 6248
rect 3516 6205 3525 6239
rect 3525 6205 3559 6239
rect 3559 6205 3568 6239
rect 3516 6196 3568 6205
rect 3884 6307 3936 6316
rect 3884 6273 3893 6307
rect 3893 6273 3927 6307
rect 3927 6273 3936 6307
rect 3884 6264 3936 6273
rect 3792 6239 3844 6248
rect 3792 6205 3801 6239
rect 3801 6205 3835 6239
rect 3835 6205 3844 6239
rect 3792 6196 3844 6205
rect 3976 6239 4028 6248
rect 3976 6205 3985 6239
rect 3985 6205 4019 6239
rect 4019 6205 4028 6239
rect 3976 6196 4028 6205
rect 4436 6375 4488 6384
rect 4436 6341 4445 6375
rect 4445 6341 4479 6375
rect 4479 6341 4488 6375
rect 4436 6332 4488 6341
rect 5540 6400 5592 6452
rect 6368 6400 6420 6452
rect 6644 6400 6696 6452
rect 6184 6332 6236 6384
rect 5540 6264 5592 6316
rect 5908 6264 5960 6316
rect 6828 6332 6880 6384
rect 7196 6400 7248 6452
rect 7380 6400 7432 6452
rect 7472 6400 7524 6452
rect 8024 6400 8076 6452
rect 8760 6400 8812 6452
rect 4436 6196 4488 6248
rect 1492 6060 1544 6112
rect 2320 6060 2372 6112
rect 3240 6060 3292 6112
rect 4344 6171 4396 6180
rect 4344 6137 4353 6171
rect 4353 6137 4387 6171
rect 4387 6137 4396 6171
rect 4344 6128 4396 6137
rect 6552 6128 6604 6180
rect 5356 6060 5408 6112
rect 6460 6060 6512 6112
rect 7012 6264 7064 6316
rect 6920 6196 6972 6248
rect 7196 6307 7248 6316
rect 7196 6273 7205 6307
rect 7205 6273 7239 6307
rect 7239 6273 7248 6307
rect 7196 6264 7248 6273
rect 7288 6196 7340 6248
rect 8024 6264 8076 6316
rect 7472 6128 7524 6180
rect 7288 6103 7340 6112
rect 7288 6069 7297 6103
rect 7297 6069 7331 6103
rect 7331 6069 7340 6103
rect 7288 6060 7340 6069
rect 7380 6060 7432 6112
rect 7840 6060 7892 6112
rect 1973 5958 2025 6010
rect 2037 5958 2089 6010
rect 2101 5958 2153 6010
rect 2165 5958 2217 6010
rect 2229 5958 2281 6010
rect 4020 5958 4072 6010
rect 4084 5958 4136 6010
rect 4148 5958 4200 6010
rect 4212 5958 4264 6010
rect 4276 5958 4328 6010
rect 6067 5958 6119 6010
rect 6131 5958 6183 6010
rect 6195 5958 6247 6010
rect 6259 5958 6311 6010
rect 6323 5958 6375 6010
rect 8114 5958 8166 6010
rect 8178 5958 8230 6010
rect 8242 5958 8294 6010
rect 8306 5958 8358 6010
rect 8370 5958 8422 6010
rect 3148 5899 3200 5908
rect 3148 5865 3157 5899
rect 3157 5865 3191 5899
rect 3191 5865 3200 5899
rect 3148 5856 3200 5865
rect 3332 5856 3384 5908
rect 3516 5856 3568 5908
rect 4344 5856 4396 5908
rect 3792 5788 3844 5840
rect 5080 5856 5132 5908
rect 5724 5856 5776 5908
rect 7104 5856 7156 5908
rect 7472 5899 7524 5908
rect 7472 5865 7481 5899
rect 7481 5865 7515 5899
rect 7515 5865 7524 5899
rect 7472 5856 7524 5865
rect 8208 5856 8260 5908
rect 2412 5720 2464 5772
rect 3240 5720 3292 5772
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 2596 5652 2648 5704
rect 3516 5763 3568 5772
rect 3516 5729 3525 5763
rect 3525 5729 3559 5763
rect 3559 5729 3568 5763
rect 3516 5720 3568 5729
rect 2504 5584 2556 5636
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 3608 5516 3660 5568
rect 4528 5720 4580 5772
rect 5264 5788 5316 5840
rect 6552 5788 6604 5840
rect 8668 5788 8720 5840
rect 5724 5763 5776 5772
rect 5724 5729 5733 5763
rect 5733 5729 5767 5763
rect 5767 5729 5776 5763
rect 5724 5720 5776 5729
rect 6736 5720 6788 5772
rect 7288 5720 7340 5772
rect 7472 5720 7524 5772
rect 8024 5720 8076 5772
rect 5080 5652 5132 5704
rect 5356 5652 5408 5704
rect 5908 5695 5960 5704
rect 5540 5584 5592 5636
rect 5908 5661 5917 5695
rect 5917 5661 5951 5695
rect 5951 5661 5960 5695
rect 5908 5652 5960 5661
rect 6276 5652 6328 5704
rect 6368 5695 6420 5704
rect 6368 5661 6377 5695
rect 6377 5661 6411 5695
rect 6411 5661 6420 5695
rect 6368 5652 6420 5661
rect 6460 5652 6512 5704
rect 6552 5652 6604 5704
rect 6828 5652 6880 5704
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 7012 5695 7064 5704
rect 7012 5661 7021 5695
rect 7021 5661 7055 5695
rect 7055 5661 7064 5695
rect 7012 5652 7064 5661
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 8760 5652 8812 5704
rect 5724 5516 5776 5568
rect 6184 5516 6236 5568
rect 7104 5516 7156 5568
rect 7932 5516 7984 5568
rect 8484 5516 8536 5568
rect 2633 5414 2685 5466
rect 2697 5414 2749 5466
rect 2761 5414 2813 5466
rect 2825 5414 2877 5466
rect 2889 5414 2941 5466
rect 4680 5414 4732 5466
rect 4744 5414 4796 5466
rect 4808 5414 4860 5466
rect 4872 5414 4924 5466
rect 4936 5414 4988 5466
rect 6727 5414 6779 5466
rect 6791 5414 6843 5466
rect 6855 5414 6907 5466
rect 6919 5414 6971 5466
rect 6983 5414 7035 5466
rect 8774 5414 8826 5466
rect 8838 5414 8890 5466
rect 8902 5414 8954 5466
rect 8966 5414 9018 5466
rect 9030 5414 9082 5466
rect 3424 5312 3476 5364
rect 3516 5312 3568 5364
rect 7196 5312 7248 5364
rect 7932 5355 7984 5364
rect 7932 5321 7941 5355
rect 7941 5321 7975 5355
rect 7975 5321 7984 5355
rect 7932 5312 7984 5321
rect 8024 5355 8076 5364
rect 8024 5321 8033 5355
rect 8033 5321 8067 5355
rect 8067 5321 8076 5355
rect 8024 5312 8076 5321
rect 8116 5312 8168 5364
rect 8208 5355 8260 5364
rect 8208 5321 8217 5355
rect 8217 5321 8251 5355
rect 8251 5321 8260 5355
rect 8208 5312 8260 5321
rect 8576 5312 8628 5364
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 3700 5244 3752 5296
rect 3056 5176 3108 5228
rect 3516 5176 3568 5228
rect 3792 5176 3844 5228
rect 4344 5219 4396 5228
rect 4344 5185 4353 5219
rect 4353 5185 4387 5219
rect 4387 5185 4396 5219
rect 4344 5176 4396 5185
rect 5172 5244 5224 5296
rect 5632 5244 5684 5296
rect 6460 5244 6512 5296
rect 7472 5244 7524 5296
rect 4068 5108 4120 5160
rect 4528 5108 4580 5160
rect 4988 5219 5040 5228
rect 4988 5185 4997 5219
rect 4997 5185 5031 5219
rect 5031 5185 5040 5219
rect 4988 5176 5040 5185
rect 5172 5108 5224 5160
rect 5816 5176 5868 5228
rect 6368 5219 6420 5228
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 6552 5219 6604 5228
rect 6552 5185 6561 5219
rect 6561 5185 6595 5219
rect 6595 5185 6604 5219
rect 6552 5176 6604 5185
rect 6828 5219 6880 5228
rect 6828 5185 6837 5219
rect 6837 5185 6871 5219
rect 6871 5185 6880 5219
rect 6828 5176 6880 5185
rect 6920 5176 6972 5228
rect 7196 5176 7248 5228
rect 7012 5108 7064 5160
rect 3424 5040 3476 5092
rect 5080 5040 5132 5092
rect 7840 5176 7892 5228
rect 8116 5219 8168 5228
rect 8116 5185 8125 5219
rect 8125 5185 8159 5219
rect 8159 5185 8168 5219
rect 8116 5176 8168 5185
rect 3608 4972 3660 5024
rect 4436 4972 4488 5024
rect 4804 4972 4856 5024
rect 5632 4972 5684 5024
rect 5816 4972 5868 5024
rect 6184 4972 6236 5024
rect 6460 5015 6512 5024
rect 6460 4981 6469 5015
rect 6469 4981 6503 5015
rect 6503 4981 6512 5015
rect 6460 4972 6512 4981
rect 6552 4972 6604 5024
rect 6736 4972 6788 5024
rect 8760 5219 8812 5228
rect 8760 5185 8769 5219
rect 8769 5185 8803 5219
rect 8803 5185 8812 5219
rect 8760 5176 8812 5185
rect 8576 5040 8628 5092
rect 7564 4972 7616 5024
rect 7840 5015 7892 5024
rect 7840 4981 7849 5015
rect 7849 4981 7883 5015
rect 7883 4981 7892 5015
rect 7840 4972 7892 4981
rect 1973 4870 2025 4922
rect 2037 4870 2089 4922
rect 2101 4870 2153 4922
rect 2165 4870 2217 4922
rect 2229 4870 2281 4922
rect 4020 4870 4072 4922
rect 4084 4870 4136 4922
rect 4148 4870 4200 4922
rect 4212 4870 4264 4922
rect 4276 4870 4328 4922
rect 6067 4870 6119 4922
rect 6131 4870 6183 4922
rect 6195 4870 6247 4922
rect 6259 4870 6311 4922
rect 6323 4870 6375 4922
rect 8114 4870 8166 4922
rect 8178 4870 8230 4922
rect 8242 4870 8294 4922
rect 8306 4870 8358 4922
rect 8370 4870 8422 4922
rect 1584 4768 1636 4820
rect 2504 4768 2556 4820
rect 4896 4768 4948 4820
rect 5264 4768 5316 4820
rect 5724 4768 5776 4820
rect 7472 4768 7524 4820
rect 8576 4768 8628 4820
rect 1584 4564 1636 4616
rect 3424 4700 3476 4752
rect 4252 4700 4304 4752
rect 6920 4700 6972 4752
rect 2412 4564 2464 4616
rect 3148 4675 3200 4684
rect 3148 4641 3157 4675
rect 3157 4641 3191 4675
rect 3191 4641 3200 4675
rect 3148 4632 3200 4641
rect 2228 4496 2280 4548
rect 3608 4564 3660 4616
rect 3700 4564 3752 4616
rect 3792 4564 3844 4616
rect 5264 4632 5316 4684
rect 5356 4675 5408 4684
rect 5356 4641 5365 4675
rect 5365 4641 5399 4675
rect 5399 4641 5408 4675
rect 5356 4632 5408 4641
rect 5632 4675 5684 4684
rect 5632 4641 5641 4675
rect 5641 4641 5675 4675
rect 5675 4641 5684 4675
rect 5632 4632 5684 4641
rect 4436 4564 4488 4616
rect 4804 4564 4856 4616
rect 4896 4564 4948 4616
rect 4988 4607 5040 4616
rect 4988 4573 4997 4607
rect 4997 4573 5031 4607
rect 5031 4573 5040 4607
rect 4988 4564 5040 4573
rect 5724 4564 5776 4616
rect 6000 4607 6052 4616
rect 6000 4573 6009 4607
rect 6009 4573 6043 4607
rect 6043 4573 6052 4607
rect 6000 4564 6052 4573
rect 6644 4607 6696 4616
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 7012 4564 7064 4616
rect 7840 4632 7892 4684
rect 7932 4632 7984 4684
rect 4160 4428 4212 4480
rect 4344 4428 4396 4480
rect 5632 4428 5684 4480
rect 6000 4428 6052 4480
rect 6736 4496 6788 4548
rect 7288 4607 7340 4616
rect 7288 4573 7297 4607
rect 7297 4573 7331 4607
rect 7331 4573 7340 4607
rect 7288 4564 7340 4573
rect 7472 4564 7524 4616
rect 8024 4607 8076 4616
rect 8024 4573 8033 4607
rect 8033 4573 8067 4607
rect 8067 4573 8076 4607
rect 8024 4564 8076 4573
rect 6276 4471 6328 4480
rect 6276 4437 6285 4471
rect 6285 4437 6319 4471
rect 6319 4437 6328 4471
rect 6276 4428 6328 4437
rect 7196 4428 7248 4480
rect 7748 4428 7800 4480
rect 8484 4607 8536 4616
rect 8484 4573 8493 4607
rect 8493 4573 8527 4607
rect 8527 4573 8536 4607
rect 8484 4564 8536 4573
rect 8300 4428 8352 4480
rect 2633 4326 2685 4378
rect 2697 4326 2749 4378
rect 2761 4326 2813 4378
rect 2825 4326 2877 4378
rect 2889 4326 2941 4378
rect 4680 4326 4732 4378
rect 4744 4326 4796 4378
rect 4808 4326 4860 4378
rect 4872 4326 4924 4378
rect 4936 4326 4988 4378
rect 6727 4326 6779 4378
rect 6791 4326 6843 4378
rect 6855 4326 6907 4378
rect 6919 4326 6971 4378
rect 6983 4326 7035 4378
rect 8774 4326 8826 4378
rect 8838 4326 8890 4378
rect 8902 4326 8954 4378
rect 8966 4326 9018 4378
rect 9030 4326 9082 4378
rect 3700 4224 3752 4276
rect 4988 4224 5040 4276
rect 5264 4224 5316 4276
rect 6460 4224 6512 4276
rect 7288 4224 7340 4276
rect 4896 4156 4948 4208
rect 5356 4156 5408 4208
rect 5448 4199 5500 4208
rect 5448 4165 5457 4199
rect 5457 4165 5491 4199
rect 5491 4165 5500 4199
rect 5448 4156 5500 4165
rect 6828 4156 6880 4208
rect 7380 4156 7432 4208
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 1676 4131 1728 4140
rect 1676 4097 1710 4131
rect 1710 4097 1728 4131
rect 1676 4088 1728 4097
rect 3240 4020 3292 4072
rect 5816 4131 5868 4140
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 7012 4088 7064 4140
rect 7472 4088 7524 4140
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 7932 4088 7984 4140
rect 5908 3952 5960 4004
rect 6644 4020 6696 4072
rect 7380 4020 7432 4072
rect 8484 4088 8536 4140
rect 8024 4020 8076 4072
rect 8300 4063 8352 4072
rect 8300 4029 8309 4063
rect 8309 4029 8343 4063
rect 8343 4029 8352 4063
rect 8300 4020 8352 4029
rect 2780 3927 2832 3936
rect 2780 3893 2789 3927
rect 2789 3893 2823 3927
rect 2823 3893 2832 3927
rect 2780 3884 2832 3893
rect 2872 3927 2924 3936
rect 2872 3893 2881 3927
rect 2881 3893 2915 3927
rect 2915 3893 2924 3927
rect 2872 3884 2924 3893
rect 3792 3884 3844 3936
rect 5264 3884 5316 3936
rect 5816 3927 5868 3936
rect 5816 3893 5825 3927
rect 5825 3893 5859 3927
rect 5859 3893 5868 3927
rect 5816 3884 5868 3893
rect 6828 3927 6880 3936
rect 6828 3893 6837 3927
rect 6837 3893 6871 3927
rect 6871 3893 6880 3927
rect 6828 3884 6880 3893
rect 7104 3884 7156 3936
rect 7932 3884 7984 3936
rect 1973 3782 2025 3834
rect 2037 3782 2089 3834
rect 2101 3782 2153 3834
rect 2165 3782 2217 3834
rect 2229 3782 2281 3834
rect 4020 3782 4072 3834
rect 4084 3782 4136 3834
rect 4148 3782 4200 3834
rect 4212 3782 4264 3834
rect 4276 3782 4328 3834
rect 6067 3782 6119 3834
rect 6131 3782 6183 3834
rect 6195 3782 6247 3834
rect 6259 3782 6311 3834
rect 6323 3782 6375 3834
rect 8114 3782 8166 3834
rect 8178 3782 8230 3834
rect 8242 3782 8294 3834
rect 8306 3782 8358 3834
rect 8370 3782 8422 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 1676 3680 1728 3732
rect 2504 3680 2556 3732
rect 5080 3680 5132 3732
rect 5264 3680 5316 3732
rect 5724 3680 5776 3732
rect 7012 3723 7064 3732
rect 7012 3689 7021 3723
rect 7021 3689 7055 3723
rect 7055 3689 7064 3723
rect 7012 3680 7064 3689
rect 7196 3680 7248 3732
rect 7380 3680 7432 3732
rect 7472 3680 7524 3732
rect 8484 3680 8536 3732
rect 3148 3612 3200 3664
rect 2412 3544 2464 3596
rect 1308 3476 1360 3528
rect 2780 3544 2832 3596
rect 3240 3544 3292 3596
rect 3792 3544 3844 3596
rect 3148 3476 3200 3528
rect 2320 3383 2372 3392
rect 2320 3349 2329 3383
rect 2329 3349 2363 3383
rect 2363 3349 2372 3383
rect 2320 3340 2372 3349
rect 2780 3383 2832 3392
rect 2780 3349 2789 3383
rect 2789 3349 2823 3383
rect 2823 3349 2832 3383
rect 2780 3340 2832 3349
rect 4160 3655 4212 3664
rect 4160 3621 4169 3655
rect 4169 3621 4203 3655
rect 4203 3621 4212 3655
rect 4160 3612 4212 3621
rect 4436 3612 4488 3664
rect 4896 3587 4948 3596
rect 4896 3553 4905 3587
rect 4905 3553 4939 3587
rect 4939 3553 4948 3587
rect 4896 3544 4948 3553
rect 4344 3519 4396 3528
rect 4344 3485 4353 3519
rect 4353 3485 4387 3519
rect 4387 3485 4396 3519
rect 4344 3476 4396 3485
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 4712 3476 4764 3528
rect 5080 3476 5132 3528
rect 5264 3451 5316 3460
rect 5264 3417 5273 3451
rect 5273 3417 5307 3451
rect 5307 3417 5316 3451
rect 5264 3408 5316 3417
rect 5540 3476 5592 3528
rect 7104 3612 7156 3664
rect 7748 3544 7800 3596
rect 6460 3476 6512 3528
rect 7380 3476 7432 3528
rect 7840 3476 7892 3528
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 7656 3408 7708 3460
rect 4712 3340 4764 3392
rect 4988 3340 5040 3392
rect 5540 3340 5592 3392
rect 2633 3238 2685 3290
rect 2697 3238 2749 3290
rect 2761 3238 2813 3290
rect 2825 3238 2877 3290
rect 2889 3238 2941 3290
rect 4680 3238 4732 3290
rect 4744 3238 4796 3290
rect 4808 3238 4860 3290
rect 4872 3238 4924 3290
rect 4936 3238 4988 3290
rect 6727 3238 6779 3290
rect 6791 3238 6843 3290
rect 6855 3238 6907 3290
rect 6919 3238 6971 3290
rect 6983 3238 7035 3290
rect 8774 3238 8826 3290
rect 8838 3238 8890 3290
rect 8902 3238 8954 3290
rect 8966 3238 9018 3290
rect 9030 3238 9082 3290
rect 2320 3136 2372 3188
rect 4252 3136 4304 3188
rect 4344 3136 4396 3188
rect 5816 3136 5868 3188
rect 7380 3136 7432 3188
rect 5080 3068 5132 3120
rect 1400 3000 1452 3052
rect 1860 3043 1912 3052
rect 1860 3009 1894 3043
rect 1894 3009 1912 3043
rect 1860 3000 1912 3009
rect 3240 3043 3292 3052
rect 3240 3009 3249 3043
rect 3249 3009 3283 3043
rect 3283 3009 3292 3043
rect 3240 3000 3292 3009
rect 3700 3000 3752 3052
rect 4252 3043 4304 3052
rect 4252 3009 4261 3043
rect 4261 3009 4295 3043
rect 4295 3009 4304 3043
rect 4252 3000 4304 3009
rect 4344 3000 4396 3052
rect 4528 3000 4580 3052
rect 5724 3043 5776 3052
rect 5724 3009 5742 3043
rect 5742 3009 5776 3043
rect 5724 3000 5776 3009
rect 5908 3000 5960 3052
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 8024 2932 8076 2984
rect 7748 2907 7800 2916
rect 7748 2873 7757 2907
rect 7757 2873 7791 2907
rect 7791 2873 7800 2907
rect 7748 2864 7800 2873
rect 3148 2796 3200 2848
rect 4620 2839 4672 2848
rect 4620 2805 4629 2839
rect 4629 2805 4663 2839
rect 4663 2805 4672 2839
rect 4620 2796 4672 2805
rect 1973 2694 2025 2746
rect 2037 2694 2089 2746
rect 2101 2694 2153 2746
rect 2165 2694 2217 2746
rect 2229 2694 2281 2746
rect 4020 2694 4072 2746
rect 4084 2694 4136 2746
rect 4148 2694 4200 2746
rect 4212 2694 4264 2746
rect 4276 2694 4328 2746
rect 6067 2694 6119 2746
rect 6131 2694 6183 2746
rect 6195 2694 6247 2746
rect 6259 2694 6311 2746
rect 6323 2694 6375 2746
rect 8114 2694 8166 2746
rect 8178 2694 8230 2746
rect 8242 2694 8294 2746
rect 8306 2694 8358 2746
rect 8370 2694 8422 2746
rect 1860 2592 1912 2644
rect 2320 2592 2372 2644
rect 2412 2635 2464 2644
rect 2412 2601 2421 2635
rect 2421 2601 2455 2635
rect 2455 2601 2464 2635
rect 2412 2592 2464 2601
rect 3516 2592 3568 2644
rect 4344 2592 4396 2644
rect 4436 2635 4488 2644
rect 4436 2601 4445 2635
rect 4445 2601 4479 2635
rect 4479 2601 4488 2635
rect 4436 2592 4488 2601
rect 5632 2592 5684 2644
rect 5724 2635 5776 2644
rect 5724 2601 5733 2635
rect 5733 2601 5767 2635
rect 5767 2601 5776 2635
rect 5724 2592 5776 2601
rect 6828 2592 6880 2644
rect 8024 2635 8076 2644
rect 8024 2601 8033 2635
rect 8033 2601 8067 2635
rect 8067 2601 8076 2635
rect 8024 2592 8076 2601
rect 3700 2524 3752 2576
rect 4528 2524 4580 2576
rect 1768 2388 1820 2440
rect 2964 2456 3016 2508
rect 3884 2456 3936 2508
rect 2780 2431 2832 2440
rect 2780 2397 2789 2431
rect 2789 2397 2823 2431
rect 2823 2397 2832 2431
rect 2780 2388 2832 2397
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 3516 2431 3568 2440
rect 3516 2397 3525 2431
rect 3525 2397 3559 2431
rect 3559 2397 3568 2431
rect 3516 2388 3568 2397
rect 3700 2388 3752 2440
rect 6644 2499 6696 2508
rect 6644 2465 6653 2499
rect 6653 2465 6687 2499
rect 6687 2465 6696 2499
rect 6644 2456 6696 2465
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 5540 2388 5592 2440
rect 2504 2252 2556 2304
rect 5172 2320 5224 2372
rect 7196 2388 7248 2440
rect 3792 2252 3844 2304
rect 2633 2150 2685 2202
rect 2697 2150 2749 2202
rect 2761 2150 2813 2202
rect 2825 2150 2877 2202
rect 2889 2150 2941 2202
rect 4680 2150 4732 2202
rect 4744 2150 4796 2202
rect 4808 2150 4860 2202
rect 4872 2150 4924 2202
rect 4936 2150 4988 2202
rect 6727 2150 6779 2202
rect 6791 2150 6843 2202
rect 6855 2150 6907 2202
rect 6919 2150 6971 2202
rect 6983 2150 7035 2202
rect 8774 2150 8826 2202
rect 8838 2150 8890 2202
rect 8902 2150 8954 2202
rect 8966 2150 9018 2202
rect 9030 2150 9082 2202
<< metal2 >>
rect 5814 11802 5870 12602
rect 1973 10364 2281 10373
rect 1973 10362 1979 10364
rect 2035 10362 2059 10364
rect 2115 10362 2139 10364
rect 2195 10362 2219 10364
rect 2275 10362 2281 10364
rect 2035 10310 2037 10362
rect 2217 10310 2219 10362
rect 1973 10308 1979 10310
rect 2035 10308 2059 10310
rect 2115 10308 2139 10310
rect 2195 10308 2219 10310
rect 2275 10308 2281 10310
rect 1973 10299 2281 10308
rect 4020 10364 4328 10373
rect 4020 10362 4026 10364
rect 4082 10362 4106 10364
rect 4162 10362 4186 10364
rect 4242 10362 4266 10364
rect 4322 10362 4328 10364
rect 4082 10310 4084 10362
rect 4264 10310 4266 10362
rect 4020 10308 4026 10310
rect 4082 10308 4106 10310
rect 4162 10308 4186 10310
rect 4242 10308 4266 10310
rect 4322 10308 4328 10310
rect 4020 10299 4328 10308
rect 5828 10266 5856 11802
rect 6067 10364 6375 10373
rect 6067 10362 6073 10364
rect 6129 10362 6153 10364
rect 6209 10362 6233 10364
rect 6289 10362 6313 10364
rect 6369 10362 6375 10364
rect 6129 10310 6131 10362
rect 6311 10310 6313 10362
rect 6067 10308 6073 10310
rect 6129 10308 6153 10310
rect 6209 10308 6233 10310
rect 6289 10308 6313 10310
rect 6369 10308 6375 10310
rect 6067 10299 6375 10308
rect 8114 10364 8422 10373
rect 8114 10362 8120 10364
rect 8176 10362 8200 10364
rect 8256 10362 8280 10364
rect 8336 10362 8360 10364
rect 8416 10362 8422 10364
rect 8176 10310 8178 10362
rect 8358 10310 8360 10362
rect 8114 10308 8120 10310
rect 8176 10308 8200 10310
rect 8256 10308 8280 10310
rect 8336 10308 8360 10310
rect 8416 10308 8422 10310
rect 8114 10299 8422 10308
rect 5816 10260 5868 10266
rect 5816 10202 5868 10208
rect 5356 10192 5408 10198
rect 5356 10134 5408 10140
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 1596 9722 1808 9738
rect 2056 9722 2084 9998
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 1584 9716 1808 9722
rect 1636 9710 1808 9716
rect 1584 9658 1636 9664
rect 1780 9674 1808 9710
rect 2044 9716 2096 9722
rect 1676 9648 1728 9654
rect 1780 9646 1900 9674
rect 2044 9658 2096 9664
rect 1676 9590 1728 9596
rect 1584 9580 1636 9586
rect 1412 9540 1584 9568
rect 1412 8974 1440 9540
rect 1584 9522 1636 9528
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1400 8968 1452 8974
rect 1596 8945 1624 9318
rect 1400 8910 1452 8916
rect 1582 8936 1638 8945
rect 1308 8492 1360 8498
rect 1308 8434 1360 8440
rect 1320 7546 1348 8434
rect 1308 7540 1360 7546
rect 1308 7482 1360 7488
rect 1412 7410 1440 8910
rect 1492 8900 1544 8906
rect 1582 8871 1638 8880
rect 1492 8842 1544 8848
rect 1504 8634 1532 8842
rect 1596 8634 1624 8871
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1492 8288 1544 8294
rect 1492 8230 1544 8236
rect 1504 8090 1532 8230
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1504 6866 1532 8026
rect 1584 8016 1636 8022
rect 1584 7958 1636 7964
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1306 6216 1362 6225
rect 1306 6151 1362 6160
rect 1320 3534 1348 6151
rect 1504 6118 1532 6802
rect 1596 6798 1624 7958
rect 1688 7750 1716 9590
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 1780 7886 1808 9454
rect 1872 8480 1900 9646
rect 1973 9276 2281 9285
rect 1973 9274 1979 9276
rect 2035 9274 2059 9276
rect 2115 9274 2139 9276
rect 2195 9274 2219 9276
rect 2275 9274 2281 9276
rect 2035 9222 2037 9274
rect 2217 9222 2219 9274
rect 1973 9220 1979 9222
rect 2035 9220 2059 9222
rect 2115 9220 2139 9222
rect 2195 9220 2219 9222
rect 2275 9220 2281 9222
rect 1973 9211 2281 9220
rect 1872 8452 1992 8480
rect 1858 8392 1914 8401
rect 1858 8327 1860 8336
rect 1912 8327 1914 8336
rect 1860 8298 1912 8304
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 1676 7744 1728 7750
rect 1728 7704 1808 7732
rect 1676 7686 1728 7692
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1688 7002 1716 7346
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1780 6798 1808 7704
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1596 6474 1624 6734
rect 1596 6446 1716 6474
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1596 6225 1624 6258
rect 1688 6254 1716 6446
rect 1872 6322 1900 8298
rect 1964 8294 1992 8452
rect 2516 8412 2544 9862
rect 2633 9820 2941 9829
rect 2633 9818 2639 9820
rect 2695 9818 2719 9820
rect 2775 9818 2799 9820
rect 2855 9818 2879 9820
rect 2935 9818 2941 9820
rect 2695 9766 2697 9818
rect 2877 9766 2879 9818
rect 2633 9764 2639 9766
rect 2695 9764 2719 9766
rect 2775 9764 2799 9766
rect 2855 9764 2879 9766
rect 2935 9764 2941 9766
rect 2633 9755 2941 9764
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2884 9178 2912 9522
rect 2976 9382 3004 9998
rect 3252 9382 3280 9998
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2976 8838 3004 9318
rect 3148 9104 3200 9110
rect 3148 9046 3200 9052
rect 3160 8974 3188 9046
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2633 8732 2941 8741
rect 2633 8730 2639 8732
rect 2695 8730 2719 8732
rect 2775 8730 2799 8732
rect 2855 8730 2879 8732
rect 2935 8730 2941 8732
rect 2695 8678 2697 8730
rect 2877 8678 2879 8730
rect 2633 8676 2639 8678
rect 2695 8676 2719 8678
rect 2775 8676 2799 8678
rect 2855 8676 2879 8678
rect 2935 8676 2941 8678
rect 2633 8667 2941 8676
rect 2976 8514 3004 8774
rect 3068 8634 3096 8910
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3056 8628 3108 8634
rect 3056 8570 3108 8576
rect 3160 8566 3188 8774
rect 2884 8486 3004 8514
rect 3148 8560 3200 8566
rect 3148 8502 3200 8508
rect 2884 8430 2912 8486
rect 2872 8424 2924 8430
rect 2424 8384 2728 8412
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 1973 8188 2281 8197
rect 1973 8186 1979 8188
rect 2035 8186 2059 8188
rect 2115 8186 2139 8188
rect 2195 8186 2219 8188
rect 2275 8186 2281 8188
rect 2035 8134 2037 8186
rect 2217 8134 2219 8186
rect 1973 8132 1979 8134
rect 2035 8132 2059 8134
rect 2115 8132 2139 8134
rect 2195 8132 2219 8134
rect 2275 8132 2281 8134
rect 1973 8123 2281 8132
rect 2318 7848 2374 7857
rect 2318 7783 2320 7792
rect 2372 7783 2374 7792
rect 2320 7754 2372 7760
rect 1973 7100 2281 7109
rect 1973 7098 1979 7100
rect 2035 7098 2059 7100
rect 2115 7098 2139 7100
rect 2195 7098 2219 7100
rect 2275 7098 2281 7100
rect 2035 7046 2037 7098
rect 2217 7046 2219 7098
rect 1973 7044 1979 7046
rect 2035 7044 2059 7046
rect 2115 7044 2139 7046
rect 2195 7044 2219 7046
rect 2275 7044 2281 7046
rect 1973 7035 2281 7044
rect 2332 6934 2360 7754
rect 2424 7478 2452 8384
rect 2700 7886 2728 8384
rect 2872 8366 2924 8372
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2792 7954 2820 8026
rect 2884 7954 2912 8366
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 2976 7993 3004 8230
rect 2962 7984 3018 7993
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2872 7948 2924 7954
rect 2962 7919 3018 7928
rect 2872 7890 2924 7896
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 2504 7812 2556 7818
rect 2504 7754 2556 7760
rect 2516 7546 2544 7754
rect 2976 7750 3004 7822
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2633 7644 2941 7653
rect 2633 7642 2639 7644
rect 2695 7642 2719 7644
rect 2775 7642 2799 7644
rect 2855 7642 2879 7644
rect 2935 7642 2941 7644
rect 2695 7590 2697 7642
rect 2877 7590 2879 7642
rect 2633 7588 2639 7590
rect 2695 7588 2719 7590
rect 2775 7588 2799 7590
rect 2855 7588 2879 7590
rect 2935 7588 2941 7590
rect 2633 7579 2941 7588
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2412 7472 2464 7478
rect 2412 7414 2464 7420
rect 2412 7268 2464 7274
rect 2412 7210 2464 7216
rect 2320 6928 2372 6934
rect 1950 6896 2006 6905
rect 2320 6870 2372 6876
rect 1950 6831 2006 6840
rect 1964 6390 1992 6831
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 2320 6792 2372 6798
rect 2320 6734 2372 6740
rect 2056 6458 2084 6734
rect 2332 6458 2360 6734
rect 2424 6730 2452 7210
rect 3068 7018 3096 8230
rect 2976 7002 3096 7018
rect 2976 6996 3108 7002
rect 2976 6990 3056 6996
rect 2412 6724 2464 6730
rect 2412 6666 2464 6672
rect 2633 6556 2941 6565
rect 2633 6554 2639 6556
rect 2695 6554 2719 6556
rect 2775 6554 2799 6556
rect 2855 6554 2879 6556
rect 2935 6554 2941 6556
rect 2695 6502 2697 6554
rect 2877 6502 2879 6554
rect 2633 6500 2639 6502
rect 2695 6500 2719 6502
rect 2775 6500 2799 6502
rect 2855 6500 2879 6502
rect 2935 6500 2941 6502
rect 2633 6491 2941 6500
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 1952 6384 2004 6390
rect 1952 6326 2004 6332
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1676 6248 1728 6254
rect 1582 6216 1638 6225
rect 1676 6190 1728 6196
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 1582 6151 1638 6160
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5234 1440 5646
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1412 4146 1440 5170
rect 1596 4826 1624 6151
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 1973 6012 2281 6021
rect 1973 6010 1979 6012
rect 2035 6010 2059 6012
rect 2115 6010 2139 6012
rect 2195 6010 2219 6012
rect 2275 6010 2281 6012
rect 2035 5958 2037 6010
rect 2217 5958 2219 6010
rect 1973 5956 1979 5958
rect 2035 5956 2059 5958
rect 2115 5956 2139 5958
rect 2195 5956 2219 5958
rect 2275 5956 2281 5958
rect 1973 5947 2281 5956
rect 1766 5264 1822 5273
rect 1766 5199 1822 5208
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1412 3058 1440 4082
rect 1596 3738 1624 4558
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 1688 3738 1716 4082
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1780 2446 1808 5199
rect 1973 4924 2281 4933
rect 1973 4922 1979 4924
rect 2035 4922 2059 4924
rect 2115 4922 2139 4924
rect 2195 4922 2219 4924
rect 2275 4922 2281 4924
rect 2035 4870 2037 4922
rect 2217 4870 2219 4922
rect 1973 4868 1979 4870
rect 2035 4868 2059 4870
rect 2115 4868 2139 4870
rect 2195 4868 2219 4870
rect 2275 4868 2281 4870
rect 1973 4859 2281 4868
rect 2228 4548 2280 4554
rect 2228 4490 2280 4496
rect 2240 4264 2268 4490
rect 2332 4434 2360 6054
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2424 4622 2452 5714
rect 2608 5710 2636 6190
rect 2596 5704 2648 5710
rect 2884 5681 2912 6394
rect 2596 5646 2648 5652
rect 2870 5672 2926 5681
rect 2504 5636 2556 5642
rect 2870 5607 2926 5616
rect 2504 5578 2556 5584
rect 2516 4826 2544 5578
rect 2633 5468 2941 5477
rect 2633 5466 2639 5468
rect 2695 5466 2719 5468
rect 2775 5466 2799 5468
rect 2855 5466 2879 5468
rect 2935 5466 2941 5468
rect 2695 5414 2697 5466
rect 2877 5414 2879 5466
rect 2633 5412 2639 5414
rect 2695 5412 2719 5414
rect 2775 5412 2799 5414
rect 2855 5412 2879 5414
rect 2935 5412 2941 5414
rect 2633 5403 2941 5412
rect 2976 5250 3004 6990
rect 3056 6938 3108 6944
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 3068 5794 3096 6802
rect 3160 6798 3188 8502
rect 3252 8362 3280 9318
rect 3436 8906 3464 9862
rect 4434 9616 4490 9625
rect 4344 9580 4396 9586
rect 4540 9602 4568 9862
rect 4680 9820 4988 9829
rect 4680 9818 4686 9820
rect 4742 9818 4766 9820
rect 4822 9818 4846 9820
rect 4902 9818 4926 9820
rect 4982 9818 4988 9820
rect 4742 9766 4744 9818
rect 4924 9766 4926 9818
rect 4680 9764 4686 9766
rect 4742 9764 4766 9766
rect 4822 9764 4846 9766
rect 4902 9764 4926 9766
rect 4982 9764 4988 9766
rect 4680 9755 4988 9764
rect 4540 9574 4660 9602
rect 4434 9551 4490 9560
rect 4344 9522 4396 9528
rect 4020 9276 4328 9285
rect 4020 9274 4026 9276
rect 4082 9274 4106 9276
rect 4162 9274 4186 9276
rect 4242 9274 4266 9276
rect 4322 9274 4328 9276
rect 4082 9222 4084 9274
rect 4264 9222 4266 9274
rect 4020 9220 4026 9222
rect 4082 9220 4106 9222
rect 4162 9220 4186 9222
rect 4242 9220 4266 9222
rect 4322 9220 4328 9222
rect 4020 9211 4328 9220
rect 3884 8968 3936 8974
rect 4160 8968 4212 8974
rect 3884 8910 3936 8916
rect 3974 8936 4030 8945
rect 3424 8900 3476 8906
rect 3424 8842 3476 8848
rect 3608 8900 3660 8906
rect 3608 8842 3660 8848
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3252 7818 3280 8298
rect 3344 8090 3372 8434
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3516 8424 3568 8430
rect 3620 8401 3648 8842
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3804 8634 3832 8774
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3896 8514 3924 8910
rect 4030 8916 4160 8922
rect 4030 8910 4212 8916
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 4030 8894 4200 8910
rect 3974 8871 4030 8880
rect 3804 8486 3924 8514
rect 3516 8366 3568 8372
rect 3606 8392 3662 8401
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3330 7984 3386 7993
rect 3436 7954 3464 8366
rect 3330 7919 3386 7928
rect 3424 7948 3476 7954
rect 3240 7812 3292 7818
rect 3240 7754 3292 7760
rect 3344 7426 3372 7919
rect 3424 7890 3476 7896
rect 3252 7398 3372 7426
rect 3252 7342 3280 7398
rect 3436 7342 3464 7890
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3252 6798 3280 7278
rect 3344 7002 3372 7278
rect 3528 7274 3556 8366
rect 3606 8327 3662 8336
rect 3608 7880 3660 7886
rect 3606 7848 3608 7857
rect 3660 7848 3662 7857
rect 3662 7806 3740 7834
rect 3606 7783 3662 7792
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3160 5914 3188 6734
rect 3252 6633 3280 6734
rect 3238 6624 3294 6633
rect 3238 6559 3294 6568
rect 3238 6488 3294 6497
rect 3238 6423 3294 6432
rect 3252 6118 3280 6423
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3344 5914 3372 6802
rect 3528 6769 3556 7210
rect 3514 6760 3570 6769
rect 3514 6695 3570 6704
rect 3516 6384 3568 6390
rect 3516 6326 3568 6332
rect 3528 6254 3556 6326
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3068 5766 3188 5794
rect 2976 5234 3096 5250
rect 2976 5228 3108 5234
rect 2976 5222 3056 5228
rect 3056 5170 3108 5176
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 3160 4690 3188 5766
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2332 4406 2544 4434
rect 2240 4236 2360 4264
rect 1973 3836 2281 3845
rect 1973 3834 1979 3836
rect 2035 3834 2059 3836
rect 2115 3834 2139 3836
rect 2195 3834 2219 3836
rect 2275 3834 2281 3836
rect 2035 3782 2037 3834
rect 2217 3782 2219 3834
rect 1973 3780 1979 3782
rect 2035 3780 2059 3782
rect 2115 3780 2139 3782
rect 2195 3780 2219 3782
rect 2275 3780 2281 3782
rect 1973 3771 2281 3780
rect 2332 3720 2360 4236
rect 2410 4040 2466 4049
rect 2410 3975 2466 3984
rect 2240 3692 2360 3720
rect 2240 3074 2268 3692
rect 2424 3602 2452 3975
rect 2516 3738 2544 4406
rect 2633 4380 2941 4389
rect 2633 4378 2639 4380
rect 2695 4378 2719 4380
rect 2775 4378 2799 4380
rect 2855 4378 2879 4380
rect 2935 4378 2941 4380
rect 2695 4326 2697 4378
rect 2877 4326 2879 4378
rect 2633 4324 2639 4326
rect 2695 4324 2719 4326
rect 2775 4324 2799 4326
rect 2855 4324 2879 4326
rect 2935 4324 2941 4326
rect 2633 4315 2941 4324
rect 3252 4162 3280 5714
rect 3330 5672 3386 5681
rect 3330 5607 3386 5616
rect 3160 4134 3280 4162
rect 2780 3936 2832 3942
rect 2780 3878 2832 3884
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2332 3194 2360 3334
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 1860 3052 1912 3058
rect 2240 3046 2360 3074
rect 1860 2994 1912 3000
rect 1872 2650 1900 2994
rect 1973 2748 2281 2757
rect 1973 2746 1979 2748
rect 2035 2746 2059 2748
rect 2115 2746 2139 2748
rect 2195 2746 2219 2748
rect 2275 2746 2281 2748
rect 2035 2694 2037 2746
rect 2217 2694 2219 2746
rect 1973 2692 1979 2694
rect 2035 2692 2059 2694
rect 2115 2692 2139 2694
rect 2195 2692 2219 2694
rect 2275 2692 2281 2694
rect 1973 2683 2281 2692
rect 2332 2650 2360 3046
rect 2424 2650 2452 3538
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 2412 2644 2464 2650
rect 2412 2586 2464 2592
rect 1768 2440 1820 2446
rect 1768 2382 1820 2388
rect 2516 2310 2544 3674
rect 2792 3602 2820 3878
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2884 3448 2912 3878
rect 3160 3670 3188 4134
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 3252 3602 3280 4014
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 3148 3528 3200 3534
rect 3148 3470 3200 3476
rect 2884 3420 3096 3448
rect 2780 3392 2832 3398
rect 2832 3352 3004 3380
rect 2780 3334 2832 3340
rect 2633 3292 2941 3301
rect 2633 3290 2639 3292
rect 2695 3290 2719 3292
rect 2775 3290 2799 3292
rect 2855 3290 2879 3292
rect 2935 3290 2941 3292
rect 2695 3238 2697 3290
rect 2877 3238 2879 3290
rect 2633 3236 2639 3238
rect 2695 3236 2719 3238
rect 2775 3236 2799 3238
rect 2855 3236 2879 3238
rect 2935 3236 2941 3238
rect 2633 3227 2941 3236
rect 2976 2774 3004 3352
rect 2792 2746 3004 2774
rect 2792 2446 2820 2746
rect 3068 2666 3096 3420
rect 3160 2854 3188 3470
rect 3252 3058 3280 3538
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 2976 2638 3096 2666
rect 2976 2514 3004 2638
rect 3160 2530 3188 2790
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 3068 2502 3188 2530
rect 3068 2446 3096 2502
rect 3252 2446 3280 2994
rect 3344 2774 3372 5607
rect 3436 5370 3464 6190
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3528 5778 3556 5850
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 3528 5370 3556 5714
rect 3620 5574 3648 7686
rect 3712 6882 3740 7806
rect 3804 7478 3832 8486
rect 4264 8362 4292 8910
rect 4356 8634 4384 9522
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3896 8090 3924 8230
rect 4020 8188 4328 8197
rect 4020 8186 4026 8188
rect 4082 8186 4106 8188
rect 4162 8186 4186 8188
rect 4242 8186 4266 8188
rect 4322 8186 4328 8188
rect 4082 8134 4084 8186
rect 4264 8134 4266 8186
rect 4020 8132 4026 8134
rect 4082 8132 4106 8134
rect 4162 8132 4186 8134
rect 4242 8132 4266 8134
rect 4322 8132 4328 8134
rect 4020 8123 4328 8132
rect 4356 8090 4384 8434
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 4020 7100 4328 7109
rect 4020 7098 4026 7100
rect 4082 7098 4106 7100
rect 4162 7098 4186 7100
rect 4242 7098 4266 7100
rect 4322 7098 4328 7100
rect 4082 7046 4084 7098
rect 4264 7046 4266 7098
rect 4020 7044 4026 7046
rect 4082 7044 4106 7046
rect 4162 7044 4186 7046
rect 4242 7044 4266 7046
rect 4322 7044 4328 7046
rect 4020 7035 4328 7044
rect 4068 6996 4120 7002
rect 4356 6984 4384 7822
rect 4068 6938 4120 6944
rect 4264 6956 4384 6984
rect 3712 6854 3832 6882
rect 3804 6848 3832 6854
rect 3804 6820 3924 6848
rect 3790 6760 3846 6769
rect 3790 6695 3846 6704
rect 3698 6624 3754 6633
rect 3698 6559 3754 6568
rect 3712 6236 3740 6559
rect 3804 6390 3832 6695
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 3896 6322 3924 6820
rect 3976 6792 4028 6798
rect 4080 6769 4108 6938
rect 4160 6792 4212 6798
rect 3976 6734 4028 6740
rect 4066 6760 4122 6769
rect 3988 6497 4016 6734
rect 4160 6734 4212 6740
rect 4066 6695 4122 6704
rect 3974 6488 4030 6497
rect 4172 6458 4200 6734
rect 3974 6423 4030 6432
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 3884 6316 3936 6322
rect 3884 6258 3936 6264
rect 3792 6248 3844 6254
rect 3712 6208 3792 6236
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3712 5302 3740 6208
rect 3976 6248 4028 6254
rect 3974 6216 3976 6225
rect 4264 6236 4292 6956
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 4028 6216 4292 6236
rect 3792 6190 3844 6196
rect 3896 6174 3974 6202
rect 4030 6208 4292 6216
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3700 5296 3752 5302
rect 3700 5238 3752 5244
rect 3804 5234 3832 5782
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3424 5092 3476 5098
rect 3424 5034 3476 5040
rect 3436 4758 3464 5034
rect 3424 4752 3476 4758
rect 3424 4694 3476 4700
rect 3344 2746 3464 2774
rect 3436 2530 3464 2746
rect 3528 2650 3556 5170
rect 3896 5148 3924 6174
rect 4356 6186 4384 6666
rect 4448 6390 4476 9551
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4540 8430 4568 9318
rect 4632 8838 4660 9574
rect 5092 9042 5120 9862
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4680 8732 4988 8741
rect 4680 8730 4686 8732
rect 4742 8730 4766 8732
rect 4822 8730 4846 8732
rect 4902 8730 4926 8732
rect 4982 8730 4988 8732
rect 4742 8678 4744 8730
rect 4924 8678 4926 8730
rect 4680 8676 4686 8678
rect 4742 8676 4766 8678
rect 4822 8676 4846 8678
rect 4902 8676 4926 8678
rect 4982 8676 4988 8678
rect 4680 8667 4988 8676
rect 5184 8634 5212 8910
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4540 7954 4568 8366
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 4540 7410 4568 7890
rect 4680 7644 4988 7653
rect 4680 7642 4686 7644
rect 4742 7642 4766 7644
rect 4822 7642 4846 7644
rect 4902 7642 4926 7644
rect 4982 7642 4988 7644
rect 4742 7590 4744 7642
rect 4924 7590 4926 7642
rect 4680 7588 4686 7590
rect 4742 7588 4766 7590
rect 4822 7588 4846 7590
rect 4902 7588 4926 7590
rect 4982 7588 4988 7590
rect 4680 7579 4988 7588
rect 5092 7528 5120 7890
rect 5000 7500 5120 7528
rect 5000 7449 5028 7500
rect 4986 7440 5042 7449
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4908 7398 4986 7426
rect 4724 6866 4752 7346
rect 4804 7268 4856 7274
rect 4804 7210 4856 7216
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4816 6798 4844 7210
rect 4908 6905 4936 7398
rect 4986 7375 5042 7384
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 4986 7032 5042 7041
rect 4986 6967 5042 6976
rect 4894 6896 4950 6905
rect 4894 6831 4950 6840
rect 4908 6798 4936 6831
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4436 6384 4488 6390
rect 4436 6326 4488 6332
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 3974 6151 4030 6160
rect 4344 6180 4396 6186
rect 4344 6122 4396 6128
rect 4020 6012 4328 6021
rect 4020 6010 4026 6012
rect 4082 6010 4106 6012
rect 4162 6010 4186 6012
rect 4242 6010 4266 6012
rect 4322 6010 4328 6012
rect 4082 5958 4084 6010
rect 4264 5958 4266 6010
rect 4020 5956 4026 5958
rect 4082 5956 4106 5958
rect 4162 5956 4186 5958
rect 4242 5956 4266 5958
rect 4322 5956 4328 5958
rect 4020 5947 4328 5956
rect 4356 5914 4384 6122
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4080 5166 4108 5646
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4068 5160 4120 5166
rect 3896 5120 4016 5148
rect 3988 5080 4016 5120
rect 4068 5102 4120 5108
rect 3804 5052 4016 5080
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3620 4622 3648 4966
rect 3804 4622 3832 5052
rect 4020 4924 4328 4933
rect 4020 4922 4026 4924
rect 4082 4922 4106 4924
rect 4162 4922 4186 4924
rect 4242 4922 4266 4924
rect 4322 4922 4328 4924
rect 4082 4870 4084 4922
rect 4264 4870 4266 4922
rect 4020 4868 4026 4870
rect 4082 4868 4106 4870
rect 4162 4868 4186 4870
rect 4242 4868 4266 4870
rect 4322 4868 4328 4870
rect 4020 4859 4328 4868
rect 4252 4752 4304 4758
rect 4252 4694 4304 4700
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3712 4282 3740 4558
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3804 3942 3832 4558
rect 4160 4480 4212 4486
rect 4264 4468 4292 4694
rect 4356 4486 4384 5170
rect 4448 5030 4476 6190
rect 4540 5778 4568 6734
rect 5000 6730 5028 6967
rect 4988 6724 5040 6730
rect 4988 6666 5040 6672
rect 4680 6556 4988 6565
rect 4680 6554 4686 6556
rect 4742 6554 4766 6556
rect 4822 6554 4846 6556
rect 4902 6554 4926 6556
rect 4982 6554 4988 6556
rect 4742 6502 4744 6554
rect 4924 6502 4926 6554
rect 4680 6500 4686 6502
rect 4742 6500 4766 6502
rect 4822 6500 4846 6502
rect 4902 6500 4926 6502
rect 4982 6500 4988 6502
rect 4680 6491 4988 6500
rect 5092 5914 5120 7346
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 4680 5468 4988 5477
rect 4680 5466 4686 5468
rect 4742 5466 4766 5468
rect 4822 5466 4846 5468
rect 4902 5466 4926 5468
rect 4982 5466 4988 5468
rect 4742 5414 4744 5466
rect 4924 5414 4926 5466
rect 4680 5412 4686 5414
rect 4742 5412 4766 5414
rect 4822 5412 4846 5414
rect 4902 5412 4926 5414
rect 4982 5412 4988 5414
rect 4680 5403 4988 5412
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4436 4616 4488 4622
rect 4434 4584 4436 4593
rect 4540 4604 4568 5102
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4816 4622 4844 4966
rect 5000 4842 5028 5170
rect 5092 5098 5120 5646
rect 5184 5302 5212 8570
rect 5276 8362 5304 9998
rect 5368 8906 5396 10134
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 6184 9988 6236 9994
rect 6184 9930 6236 9936
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 6196 9722 6224 9930
rect 6727 9820 7035 9829
rect 6727 9818 6733 9820
rect 6789 9818 6813 9820
rect 6869 9818 6893 9820
rect 6949 9818 6973 9820
rect 7029 9818 7035 9820
rect 6789 9766 6791 9818
rect 6971 9766 6973 9818
rect 6727 9764 6733 9766
rect 6789 9764 6813 9766
rect 6869 9764 6893 9766
rect 6949 9764 6973 9766
rect 7029 9764 7035 9766
rect 6727 9755 7035 9764
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 5724 9648 5776 9654
rect 5724 9590 5776 9596
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5460 9178 5488 9522
rect 5540 9376 5592 9382
rect 5592 9336 5672 9364
rect 5540 9318 5592 9324
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5644 8974 5672 9336
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5552 8498 5580 8842
rect 5736 8634 5764 9590
rect 6196 9586 6224 9658
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6067 9276 6375 9285
rect 6067 9274 6073 9276
rect 6129 9274 6153 9276
rect 6209 9274 6233 9276
rect 6289 9274 6313 9276
rect 6369 9274 6375 9276
rect 6129 9222 6131 9274
rect 6311 9222 6313 9274
rect 6067 9220 6073 9222
rect 6129 9220 6153 9222
rect 6209 9220 6233 9222
rect 6289 9220 6313 9222
rect 6369 9220 6375 9222
rect 6067 9211 6375 9220
rect 6000 9172 6052 9178
rect 6472 9166 6868 9194
rect 6472 9160 6500 9166
rect 6000 9114 6052 9120
rect 6380 9132 6500 9160
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5828 8514 5856 8774
rect 5920 8566 5948 8774
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5736 8486 5856 8514
rect 5908 8560 5960 8566
rect 5908 8502 5960 8508
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5368 7886 5396 8230
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5354 7576 5410 7585
rect 5354 7511 5356 7520
rect 5408 7511 5410 7520
rect 5356 7482 5408 7488
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5276 6934 5304 7346
rect 5368 7002 5396 7346
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5264 6928 5316 6934
rect 5264 6870 5316 6876
rect 5368 6746 5396 6938
rect 5276 6718 5396 6746
rect 5276 5846 5304 6718
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5368 6118 5396 6598
rect 5460 6440 5488 8434
rect 5552 7936 5580 8434
rect 5736 8090 5764 8486
rect 6012 8412 6040 9114
rect 6184 8968 6236 8974
rect 6182 8936 6184 8945
rect 6276 8968 6328 8974
rect 6236 8936 6238 8945
rect 6276 8910 6328 8916
rect 6182 8871 6238 8880
rect 5920 8384 6040 8412
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5920 8022 5948 8384
rect 6288 8294 6316 8910
rect 6380 8498 6408 9132
rect 6840 8974 6868 9166
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6644 8968 6696 8974
rect 6564 8928 6644 8956
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6067 8188 6375 8197
rect 6067 8186 6073 8188
rect 6129 8186 6153 8188
rect 6209 8186 6233 8188
rect 6289 8186 6313 8188
rect 6369 8186 6375 8188
rect 6129 8134 6131 8186
rect 6311 8134 6313 8186
rect 6067 8132 6073 8134
rect 6129 8132 6153 8134
rect 6209 8132 6233 8134
rect 6289 8132 6313 8134
rect 6369 8132 6375 8134
rect 6067 8123 6375 8132
rect 5908 8016 5960 8022
rect 5908 7958 5960 7964
rect 6184 8016 6236 8022
rect 6184 7958 6236 7964
rect 5552 7908 5672 7936
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5552 7002 5580 7754
rect 5644 7546 5672 7908
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5552 6798 5580 6938
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5540 6452 5592 6458
rect 5460 6412 5540 6440
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5264 5840 5316 5846
rect 5264 5782 5316 5788
rect 5356 5704 5408 5710
rect 5354 5672 5356 5681
rect 5408 5672 5410 5681
rect 5354 5607 5410 5616
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 4908 4826 5028 4842
rect 4896 4820 5028 4826
rect 4948 4814 5028 4820
rect 4896 4762 4948 4768
rect 5092 4706 5120 5034
rect 5000 4678 5120 4706
rect 5000 4622 5028 4678
rect 4488 4584 4568 4604
rect 4490 4576 4568 4584
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 4434 4519 4490 4528
rect 4212 4440 4292 4468
rect 4344 4480 4396 4486
rect 4160 4422 4212 4428
rect 4908 4468 4936 4558
rect 4908 4440 5120 4468
rect 4344 4422 4396 4428
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3804 3602 3832 3878
rect 4020 3836 4328 3845
rect 4020 3834 4026 3836
rect 4082 3834 4106 3836
rect 4162 3834 4186 3836
rect 4242 3834 4266 3836
rect 4322 3834 4328 3836
rect 4082 3782 4084 3834
rect 4264 3782 4266 3834
rect 4020 3780 4026 3782
rect 4082 3780 4106 3782
rect 4162 3780 4186 3782
rect 4242 3780 4266 3782
rect 4322 3780 4328 3782
rect 4020 3771 4328 3780
rect 4160 3664 4212 3670
rect 4356 3618 4384 4422
rect 4680 4380 4988 4389
rect 4680 4378 4686 4380
rect 4742 4378 4766 4380
rect 4822 4378 4846 4380
rect 4902 4378 4926 4380
rect 4982 4378 4988 4380
rect 4742 4326 4744 4378
rect 4924 4326 4926 4378
rect 4680 4324 4686 4326
rect 4742 4324 4766 4326
rect 4822 4324 4846 4326
rect 4902 4324 4926 4326
rect 4982 4324 4988 4326
rect 4680 4315 4988 4324
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 4896 4208 4948 4214
rect 4896 4150 4948 4156
rect 4160 3606 4212 3612
rect 3792 3596 3844 3602
rect 3792 3538 3844 3544
rect 4172 3074 4200 3606
rect 4264 3590 4384 3618
rect 4436 3664 4488 3670
rect 4436 3606 4488 3612
rect 4264 3194 4292 3590
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 4356 3194 4384 3470
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4344 3188 4396 3194
rect 4344 3130 4396 3136
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3804 3046 4200 3074
rect 4252 3052 4304 3058
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3712 2582 3740 2994
rect 3700 2576 3752 2582
rect 3436 2502 3556 2530
rect 3700 2518 3752 2524
rect 3528 2446 3556 2502
rect 3712 2446 3740 2518
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3700 2440 3752 2446
rect 3700 2382 3752 2388
rect 3804 2310 3832 3046
rect 4252 2994 4304 3000
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4264 2938 4292 2994
rect 3896 2910 4292 2938
rect 3896 2514 3924 2910
rect 4020 2748 4328 2757
rect 4020 2746 4026 2748
rect 4082 2746 4106 2748
rect 4162 2746 4186 2748
rect 4242 2746 4266 2748
rect 4322 2746 4328 2748
rect 4082 2694 4084 2746
rect 4264 2694 4266 2746
rect 4020 2692 4026 2694
rect 4082 2692 4106 2694
rect 4162 2692 4186 2694
rect 4242 2692 4266 2694
rect 4322 2692 4328 2694
rect 4020 2683 4328 2692
rect 4356 2650 4384 2994
rect 4448 2650 4476 3606
rect 4908 3602 4936 4150
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 4528 3528 4580 3534
rect 4712 3528 4764 3534
rect 4528 3470 4580 3476
rect 4710 3496 4712 3505
rect 4764 3496 4766 3505
rect 4540 3058 4568 3470
rect 4710 3431 4766 3440
rect 4724 3398 4752 3431
rect 5000 3398 5028 4218
rect 5092 3738 5120 4440
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5080 3528 5132 3534
rect 5184 3482 5212 5102
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5276 4690 5304 4762
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5276 4282 5304 4626
rect 5264 4276 5316 4282
rect 5264 4218 5316 4224
rect 5368 4214 5396 4626
rect 5460 4214 5488 6412
rect 5540 6394 5592 6400
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5552 5642 5580 6258
rect 5644 5760 5672 7482
rect 5736 5914 5764 7754
rect 5828 7750 5856 7822
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5724 5772 5776 5778
rect 5644 5732 5724 5760
rect 5724 5714 5776 5720
rect 5540 5636 5592 5642
rect 5540 5578 5592 5584
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5644 5030 5672 5238
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5644 4690 5672 4966
rect 5736 4826 5764 5510
rect 5828 5234 5856 7686
rect 5920 6322 5948 7822
rect 5998 7440 6054 7449
rect 6196 7410 6224 7958
rect 6564 7954 6592 8928
rect 6644 8910 6696 8916
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6932 8820 6960 9114
rect 7116 8922 7144 9930
rect 7208 9586 7236 9998
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7300 9178 7328 10066
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7116 8894 7236 8922
rect 6656 8792 6960 8820
rect 7104 8832 7156 8838
rect 6656 8498 6684 8792
rect 7104 8774 7156 8780
rect 6727 8732 7035 8741
rect 6727 8730 6733 8732
rect 6789 8730 6813 8732
rect 6869 8730 6893 8732
rect 6949 8730 6973 8732
rect 7029 8730 7035 8732
rect 6789 8678 6791 8730
rect 6971 8678 6973 8730
rect 6727 8676 6733 8678
rect 6789 8676 6813 8678
rect 6869 8676 6893 8678
rect 6949 8676 6973 8678
rect 7029 8676 7035 8678
rect 6727 8667 7035 8676
rect 7116 8634 7144 8774
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6288 7410 6316 7686
rect 6656 7426 6684 8298
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6748 7886 6776 8230
rect 7208 8090 7236 8894
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7300 8090 7328 8434
rect 7392 8430 7420 9522
rect 7484 9178 7512 9930
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7576 8945 7604 9998
rect 7668 9654 7696 10134
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7852 9042 7880 9862
rect 8036 9382 8064 9930
rect 8774 9820 9082 9829
rect 8774 9818 8780 9820
rect 8836 9818 8860 9820
rect 8916 9818 8940 9820
rect 8996 9818 9020 9820
rect 9076 9818 9082 9820
rect 8836 9766 8838 9818
rect 9018 9766 9020 9818
rect 8774 9764 8780 9766
rect 8836 9764 8860 9766
rect 8916 9764 8940 9766
rect 8996 9764 9020 9766
rect 9076 9764 9082 9766
rect 8774 9755 9082 9764
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 7840 9036 7892 9042
rect 7840 8978 7892 8984
rect 7656 8968 7708 8974
rect 7562 8936 7618 8945
rect 7656 8910 7708 8916
rect 7562 8871 7618 8880
rect 7472 8628 7524 8634
rect 7472 8570 7524 8576
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 6932 7886 6960 7958
rect 7208 7886 7236 8026
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6920 7880 6972 7886
rect 7196 7880 7248 7886
rect 6972 7840 7144 7868
rect 6920 7822 6972 7828
rect 6748 7750 6776 7822
rect 6736 7744 6788 7750
rect 7116 7732 7144 7840
rect 7196 7822 7248 7828
rect 7116 7704 7236 7732
rect 6736 7686 6788 7692
rect 6727 7644 7035 7653
rect 6727 7642 6733 7644
rect 6789 7642 6813 7644
rect 6869 7642 6893 7644
rect 6949 7642 6973 7644
rect 7029 7642 7035 7644
rect 6789 7590 6791 7642
rect 6971 7590 6973 7642
rect 6727 7588 6733 7590
rect 6789 7588 6813 7590
rect 6869 7588 6893 7590
rect 6949 7588 6973 7590
rect 7029 7588 7035 7590
rect 6727 7579 7035 7588
rect 5998 7375 6054 7384
rect 6184 7404 6236 7410
rect 6012 7274 6040 7375
rect 6184 7346 6236 7352
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6472 7398 6684 7426
rect 6736 7404 6788 7410
rect 6000 7268 6052 7274
rect 6000 7210 6052 7216
rect 6276 7200 6328 7206
rect 6472 7188 6500 7398
rect 6736 7346 6788 7352
rect 6328 7160 6500 7188
rect 6276 7142 6328 7148
rect 6067 7100 6375 7109
rect 6067 7098 6073 7100
rect 6129 7098 6153 7100
rect 6209 7098 6233 7100
rect 6289 7098 6313 7100
rect 6369 7098 6375 7100
rect 6129 7046 6131 7098
rect 6311 7046 6313 7098
rect 6067 7044 6073 7046
rect 6129 7044 6153 7046
rect 6209 7044 6233 7046
rect 6289 7044 6313 7046
rect 6369 7044 6375 7046
rect 6067 7035 6375 7044
rect 6182 6896 6238 6905
rect 6182 6831 6238 6840
rect 6276 6860 6328 6866
rect 6196 6390 6224 6831
rect 6276 6802 6328 6808
rect 6184 6384 6236 6390
rect 6184 6326 6236 6332
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 6288 6100 6316 6802
rect 6368 6724 6420 6730
rect 6368 6666 6420 6672
rect 6380 6458 6408 6666
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6366 6216 6422 6225
rect 6472 6202 6500 7160
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6564 6338 6592 7142
rect 6656 6458 6684 7142
rect 6748 6934 6776 7346
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6840 7002 6868 7142
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6828 6792 6880 6798
rect 6826 6760 6828 6769
rect 7104 6792 7156 6798
rect 6880 6760 6882 6769
rect 7104 6734 7156 6740
rect 6826 6695 6882 6704
rect 6727 6556 7035 6565
rect 6727 6554 6733 6556
rect 6789 6554 6813 6556
rect 6869 6554 6893 6556
rect 6949 6554 6973 6556
rect 7029 6554 7035 6556
rect 6789 6502 6791 6554
rect 6971 6502 6973 6554
rect 6727 6500 6733 6502
rect 6789 6500 6813 6502
rect 6869 6500 6893 6502
rect 6949 6500 6973 6502
rect 7029 6500 7035 6502
rect 6727 6491 7035 6500
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6828 6384 6880 6390
rect 6564 6310 6684 6338
rect 6828 6326 6880 6332
rect 6422 6174 6500 6202
rect 6552 6180 6604 6186
rect 6366 6151 6422 6160
rect 6552 6122 6604 6128
rect 6460 6112 6512 6118
rect 6288 6072 6460 6100
rect 6460 6054 6512 6060
rect 6067 6012 6375 6021
rect 6067 6010 6073 6012
rect 6129 6010 6153 6012
rect 6209 6010 6233 6012
rect 6289 6010 6313 6012
rect 6369 6010 6375 6012
rect 6129 5958 6131 6010
rect 6311 5958 6313 6010
rect 6067 5956 6073 5958
rect 6129 5956 6153 5958
rect 6209 5956 6233 5958
rect 6289 5956 6313 5958
rect 6369 5956 6375 5958
rect 6067 5947 6375 5956
rect 6472 5896 6500 6054
rect 6380 5868 6500 5896
rect 6380 5710 6408 5868
rect 6564 5846 6592 6122
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5816 5024 5868 5030
rect 5816 4966 5868 4972
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5724 4616 5776 4622
rect 5722 4584 5724 4593
rect 5776 4584 5778 4593
rect 5722 4519 5778 4528
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 5448 4208 5500 4214
rect 5448 4150 5500 4156
rect 5644 4049 5672 4422
rect 5828 4146 5856 4966
rect 5920 4842 5948 5646
rect 6184 5568 6236 5574
rect 6184 5510 6236 5516
rect 6196 5030 6224 5510
rect 6288 5273 6316 5646
rect 6274 5264 6330 5273
rect 6380 5234 6408 5646
rect 6472 5302 6500 5646
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6564 5234 6592 5646
rect 6274 5199 6330 5208
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6552 5024 6604 5030
rect 6656 5012 6684 6310
rect 6734 6216 6790 6225
rect 6734 6151 6790 6160
rect 6748 5778 6776 6151
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6840 5710 6868 6326
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6932 5710 6960 6190
rect 7024 5710 7052 6258
rect 7116 5914 7144 6734
rect 7208 6458 7236 7704
rect 7286 7440 7342 7449
rect 7286 7375 7288 7384
rect 7340 7375 7342 7384
rect 7288 7346 7340 7352
rect 7392 6866 7420 8366
rect 7484 8090 7512 8570
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7484 7426 7512 8026
rect 7576 7970 7604 8871
rect 7668 8634 7696 8910
rect 7852 8838 7880 8978
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7668 8090 7696 8434
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 8036 8022 8064 9318
rect 8114 9276 8422 9285
rect 8114 9274 8120 9276
rect 8176 9274 8200 9276
rect 8256 9274 8280 9276
rect 8336 9274 8360 9276
rect 8416 9274 8422 9276
rect 8176 9222 8178 9274
rect 8358 9222 8360 9274
rect 8114 9220 8120 9222
rect 8176 9220 8200 9222
rect 8256 9220 8280 9222
rect 8336 9220 8360 9222
rect 8416 9220 8422 9222
rect 8114 9211 8422 9220
rect 8774 8732 9082 8741
rect 8774 8730 8780 8732
rect 8836 8730 8860 8732
rect 8916 8730 8940 8732
rect 8996 8730 9020 8732
rect 9076 8730 9082 8732
rect 8836 8678 8838 8730
rect 9018 8678 9020 8730
rect 8774 8676 8780 8678
rect 8836 8676 8860 8678
rect 8916 8676 8940 8678
rect 8996 8676 9020 8678
rect 9076 8676 9082 8678
rect 8774 8667 9082 8676
rect 8114 8188 8422 8197
rect 8114 8186 8120 8188
rect 8176 8186 8200 8188
rect 8256 8186 8280 8188
rect 8336 8186 8360 8188
rect 8416 8186 8422 8188
rect 8176 8134 8178 8186
rect 8358 8134 8360 8186
rect 8114 8132 8120 8134
rect 8176 8132 8200 8134
rect 8256 8132 8280 8134
rect 8336 8132 8360 8134
rect 8416 8132 8422 8134
rect 8114 8123 8422 8132
rect 8024 8016 8076 8022
rect 7576 7942 7788 7970
rect 8024 7958 8076 7964
rect 7576 7546 7604 7942
rect 7760 7886 7788 7942
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7564 7540 7616 7546
rect 7564 7482 7616 7488
rect 7484 7398 7604 7426
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7392 6458 7420 6802
rect 7484 6798 7512 7142
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7484 6458 7512 6598
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 6727 5468 7035 5477
rect 6727 5466 6733 5468
rect 6789 5466 6813 5468
rect 6869 5466 6893 5468
rect 6949 5466 6973 5468
rect 7029 5466 7035 5468
rect 6789 5414 6791 5466
rect 6971 5414 6973 5466
rect 6727 5412 6733 5414
rect 6789 5412 6813 5414
rect 6869 5412 6893 5414
rect 6949 5412 6973 5414
rect 7029 5412 7035 5414
rect 6727 5403 7035 5412
rect 7116 5250 7144 5510
rect 7208 5370 7236 6258
rect 7288 6248 7340 6254
rect 7340 6196 7420 6202
rect 7288 6190 7420 6196
rect 7300 6174 7420 6190
rect 7392 6118 7420 6174
rect 7472 6180 7524 6186
rect 7472 6122 7524 6128
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7300 5896 7328 6054
rect 7484 5914 7512 6122
rect 7472 5908 7524 5914
rect 7300 5868 7420 5896
rect 7288 5772 7340 5778
rect 7392 5760 7420 5868
rect 7472 5850 7524 5856
rect 7472 5772 7524 5778
rect 7392 5732 7472 5760
rect 7288 5714 7340 5720
rect 7472 5714 7524 5720
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 7024 5222 7144 5250
rect 7196 5228 7248 5234
rect 6736 5024 6788 5030
rect 6656 4984 6736 5012
rect 6552 4966 6604 4972
rect 6736 4966 6788 4972
rect 6067 4924 6375 4933
rect 6067 4922 6073 4924
rect 6129 4922 6153 4924
rect 6209 4922 6233 4924
rect 6289 4922 6313 4924
rect 6369 4922 6375 4924
rect 6129 4870 6131 4922
rect 6311 4870 6313 4922
rect 6067 4868 6073 4870
rect 6129 4868 6153 4870
rect 6209 4868 6233 4870
rect 6289 4868 6313 4870
rect 6369 4868 6375 4870
rect 6067 4859 6375 4868
rect 5920 4814 6040 4842
rect 6012 4622 6040 4814
rect 6274 4720 6330 4729
rect 6274 4655 6330 4664
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6012 4486 6040 4558
rect 6288 4486 6316 4655
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 6472 4282 6500 4966
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5630 4040 5686 4049
rect 5828 4026 5856 4082
rect 5630 3975 5686 3984
rect 5736 3998 5856 4026
rect 5908 4004 5960 4010
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5276 3738 5304 3878
rect 5736 3738 5764 3998
rect 5908 3946 5960 3952
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5264 3732 5316 3738
rect 5724 3732 5776 3738
rect 5264 3674 5316 3680
rect 5644 3692 5724 3720
rect 5540 3528 5592 3534
rect 5132 3476 5212 3482
rect 5080 3470 5212 3476
rect 5092 3454 5212 3470
rect 5538 3496 5540 3505
rect 5592 3496 5594 3505
rect 5264 3460 5316 3466
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4680 3292 4988 3301
rect 4680 3290 4686 3292
rect 4742 3290 4766 3292
rect 4822 3290 4846 3292
rect 4902 3290 4926 3292
rect 4982 3290 4988 3292
rect 4742 3238 4744 3290
rect 4924 3238 4926 3290
rect 4680 3236 4686 3238
rect 4742 3236 4766 3238
rect 4822 3236 4846 3238
rect 4902 3236 4926 3238
rect 4982 3236 4988 3238
rect 4680 3227 4988 3236
rect 5092 3126 5120 3454
rect 5538 3431 5594 3440
rect 5264 3402 5316 3408
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4620 2848 4672 2854
rect 4540 2796 4620 2802
rect 4540 2790 4672 2796
rect 4540 2774 4660 2790
rect 5276 2774 5304 3402
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4540 2582 4568 2774
rect 5276 2746 5488 2774
rect 4528 2576 4580 2582
rect 4528 2518 4580 2524
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 5460 2446 5488 2746
rect 5552 2446 5580 3334
rect 5644 2650 5672 3692
rect 5724 3674 5776 3680
rect 5828 3194 5856 3878
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 5920 3058 5948 3946
rect 6067 3836 6375 3845
rect 6067 3834 6073 3836
rect 6129 3834 6153 3836
rect 6209 3834 6233 3836
rect 6289 3834 6313 3836
rect 6369 3834 6375 3836
rect 6129 3782 6131 3834
rect 6311 3782 6313 3834
rect 6067 3780 6073 3782
rect 6129 3780 6153 3782
rect 6209 3780 6233 3782
rect 6289 3780 6313 3782
rect 6369 3780 6375 3782
rect 6067 3771 6375 3780
rect 6472 3534 6500 4218
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 5736 2650 5764 2994
rect 6380 2938 6408 2994
rect 6380 2910 6500 2938
rect 6067 2748 6375 2757
rect 6067 2746 6073 2748
rect 6129 2746 6153 2748
rect 6209 2746 6233 2748
rect 6289 2746 6313 2748
rect 6369 2746 6375 2748
rect 6129 2694 6131 2746
rect 6311 2694 6313 2746
rect 6067 2692 6073 2694
rect 6129 2692 6153 2694
rect 6209 2692 6233 2694
rect 6289 2692 6313 2694
rect 6369 2692 6375 2694
rect 6067 2683 6375 2692
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5724 2644 5776 2650
rect 6472 2632 6500 2910
rect 6564 2774 6592 4966
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6656 4078 6684 4558
rect 6748 4554 6776 4966
rect 6736 4548 6788 4554
rect 6736 4490 6788 4496
rect 6840 4468 6868 5170
rect 6932 4758 6960 5170
rect 7024 5166 7052 5222
rect 7300 5216 7328 5714
rect 7470 5672 7526 5681
rect 7576 5658 7604 7398
rect 7656 7268 7708 7274
rect 7656 7210 7708 7216
rect 7668 6798 7696 7210
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7526 5630 7604 5658
rect 7470 5607 7526 5616
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 7248 5188 7328 5216
rect 7196 5170 7248 5176
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 7024 4622 7052 5102
rect 7484 4826 7512 5238
rect 7760 5216 7788 7686
rect 7944 7546 7972 7686
rect 8312 7546 8340 7822
rect 8774 7644 9082 7653
rect 8774 7642 8780 7644
rect 8836 7642 8860 7644
rect 8916 7642 8940 7644
rect 8996 7642 9020 7644
rect 9076 7642 9082 7644
rect 8836 7590 8838 7642
rect 9018 7590 9020 7642
rect 8774 7588 8780 7590
rect 8836 7588 8860 7590
rect 8916 7588 8940 7590
rect 8996 7588 9020 7590
rect 9076 7588 9082 7590
rect 8774 7579 9082 7588
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 8760 7336 8812 7342
rect 8760 7278 8812 7284
rect 8036 6458 8064 7278
rect 8114 7100 8422 7109
rect 8114 7098 8120 7100
rect 8176 7098 8200 7100
rect 8256 7098 8280 7100
rect 8336 7098 8360 7100
rect 8416 7098 8422 7100
rect 8176 7046 8178 7098
rect 8358 7046 8360 7098
rect 8114 7044 8120 7046
rect 8176 7044 8200 7046
rect 8256 7044 8280 7046
rect 8336 7044 8360 7046
rect 8416 7044 8422 7046
rect 8114 7035 8422 7044
rect 8772 7002 8800 7278
rect 8760 6996 8812 7002
rect 8760 6938 8812 6944
rect 8772 6746 8800 6938
rect 8576 6724 8628 6730
rect 8576 6666 8628 6672
rect 8680 6718 8800 6746
rect 8024 6452 8076 6458
rect 7852 6412 8024 6440
rect 7852 6118 7880 6412
rect 8024 6394 8076 6400
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 5234 7880 6054
rect 8036 5778 8064 6258
rect 8114 6012 8422 6021
rect 8114 6010 8120 6012
rect 8176 6010 8200 6012
rect 8256 6010 8280 6012
rect 8336 6010 8360 6012
rect 8416 6010 8422 6012
rect 8176 5958 8178 6010
rect 8358 5958 8360 6010
rect 8114 5956 8120 5958
rect 8176 5956 8200 5958
rect 8256 5956 8280 5958
rect 8336 5956 8360 5958
rect 8416 5956 8422 5958
rect 8114 5947 8422 5956
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7944 5370 7972 5510
rect 8036 5370 8064 5714
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8128 5370 8156 5646
rect 8220 5370 8248 5850
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8036 5250 8064 5306
rect 7668 5188 7788 5216
rect 7840 5228 7892 5234
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7484 4622 7512 4762
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7288 4616 7340 4622
rect 7472 4616 7524 4622
rect 7288 4558 7340 4564
rect 7392 4576 7472 4604
rect 7196 4480 7248 4486
rect 6840 4440 7144 4468
rect 6727 4380 7035 4389
rect 6727 4378 6733 4380
rect 6789 4378 6813 4380
rect 6869 4378 6893 4380
rect 6949 4378 6973 4380
rect 7029 4378 7035 4380
rect 6789 4326 6791 4378
rect 6971 4326 6973 4378
rect 6727 4324 6733 4326
rect 6789 4324 6813 4326
rect 6869 4324 6893 4326
rect 6949 4324 6973 4326
rect 7029 4324 7035 4326
rect 6727 4315 7035 4324
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6840 3942 6868 4150
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 7024 3738 7052 4082
rect 7116 3942 7144 4440
rect 7196 4422 7248 4428
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7208 3738 7236 4422
rect 7300 4282 7328 4558
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7392 4214 7420 4576
rect 7472 4558 7524 4564
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7576 4146 7604 4966
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7392 3738 7420 4014
rect 7484 3738 7512 4082
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7196 3732 7248 3738
rect 7196 3674 7248 3680
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7472 3732 7524 3738
rect 7472 3674 7524 3680
rect 7104 3664 7156 3670
rect 7104 3606 7156 3612
rect 6727 3292 7035 3301
rect 6727 3290 6733 3292
rect 6789 3290 6813 3292
rect 6869 3290 6893 3292
rect 6949 3290 6973 3292
rect 7029 3290 7035 3292
rect 6789 3238 6791 3290
rect 6971 3238 6973 3290
rect 6727 3236 6733 3238
rect 6789 3236 6813 3238
rect 6869 3236 6893 3238
rect 6949 3236 6973 3238
rect 7029 3236 7035 3238
rect 6727 3227 7035 3236
rect 7116 2774 7144 3606
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7392 3194 7420 3470
rect 7668 3466 7696 5188
rect 7840 5170 7892 5176
rect 7944 5222 8064 5250
rect 8116 5228 8168 5234
rect 7852 5114 7880 5170
rect 7760 5086 7880 5114
rect 7760 4486 7788 5086
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7852 4690 7880 4966
rect 7944 4690 7972 5222
rect 8116 5170 8168 5176
rect 8128 5114 8156 5170
rect 8036 5086 8156 5114
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 7932 4684 7984 4690
rect 7932 4626 7984 4632
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 7760 3720 7788 4422
rect 7944 4146 7972 4626
rect 8036 4622 8064 5086
rect 8114 4924 8422 4933
rect 8114 4922 8120 4924
rect 8176 4922 8200 4924
rect 8256 4922 8280 4924
rect 8336 4922 8360 4924
rect 8416 4922 8422 4924
rect 8176 4870 8178 4922
rect 8358 4870 8360 4922
rect 8114 4868 8120 4870
rect 8176 4868 8200 4870
rect 8256 4868 8280 4870
rect 8336 4868 8360 4870
rect 8416 4868 8422 4870
rect 8114 4859 8422 4868
rect 8496 4622 8524 5510
rect 8588 5370 8616 6666
rect 8680 5846 8708 6718
rect 8774 6556 9082 6565
rect 8774 6554 8780 6556
rect 8836 6554 8860 6556
rect 8916 6554 8940 6556
rect 8996 6554 9020 6556
rect 9076 6554 9082 6556
rect 8836 6502 8838 6554
rect 9018 6502 9020 6554
rect 8774 6500 8780 6502
rect 8836 6500 8860 6502
rect 8916 6500 8940 6502
rect 8996 6500 9020 6502
rect 9076 6500 9082 6502
rect 8774 6491 9082 6500
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8668 5840 8720 5846
rect 8668 5782 8720 5788
rect 8772 5710 8800 6394
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8774 5468 9082 5477
rect 8774 5466 8780 5468
rect 8836 5466 8860 5468
rect 8916 5466 8940 5468
rect 8996 5466 9020 5468
rect 9076 5466 9082 5468
rect 8836 5414 8838 5466
rect 9018 5414 9020 5466
rect 8774 5412 8780 5414
rect 8836 5412 8860 5414
rect 8916 5412 8940 5414
rect 8996 5412 9020 5414
rect 9076 5412 9082 5414
rect 8774 5403 9082 5412
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8758 5264 8814 5273
rect 8758 5199 8760 5208
rect 8812 5199 8814 5208
rect 8760 5170 8812 5176
rect 8576 5092 8628 5098
rect 8576 5034 8628 5040
rect 8588 4826 8616 5034
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 8036 4078 8064 4558
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8312 4078 8340 4422
rect 8496 4146 8524 4558
rect 8774 4380 9082 4389
rect 8774 4378 8780 4380
rect 8836 4378 8860 4380
rect 8916 4378 8940 4380
rect 8996 4378 9020 4380
rect 9076 4378 9082 4380
rect 8836 4326 8838 4378
rect 9018 4326 9020 4378
rect 8774 4324 8780 4326
rect 8836 4324 8860 4326
rect 8916 4324 8940 4326
rect 8996 4324 9020 4326
rect 9076 4324 9082 4326
rect 8774 4315 9082 4324
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7760 3692 7880 3720
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7760 2922 7788 3538
rect 7852 3534 7880 3692
rect 7944 3534 7972 3878
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 8036 2990 8064 4014
rect 8114 3836 8422 3845
rect 8114 3834 8120 3836
rect 8176 3834 8200 3836
rect 8256 3834 8280 3836
rect 8336 3834 8360 3836
rect 8416 3834 8422 3836
rect 8176 3782 8178 3834
rect 8358 3782 8360 3834
rect 8114 3780 8120 3782
rect 8176 3780 8200 3782
rect 8256 3780 8280 3782
rect 8336 3780 8360 3782
rect 8416 3780 8422 3782
rect 8114 3771 8422 3780
rect 8496 3738 8524 4082
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8774 3292 9082 3301
rect 8774 3290 8780 3292
rect 8836 3290 8860 3292
rect 8916 3290 8940 3292
rect 8996 3290 9020 3292
rect 9076 3290 9082 3292
rect 8836 3238 8838 3290
rect 9018 3238 9020 3290
rect 8774 3236 8780 3238
rect 8836 3236 8860 3238
rect 8916 3236 8940 3238
rect 8996 3236 9020 3238
rect 9076 3236 9082 3238
rect 8774 3227 9082 3236
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 6564 2746 6868 2774
rect 7116 2746 7236 2774
rect 6840 2650 6868 2746
rect 6828 2644 6880 2650
rect 6472 2604 6684 2632
rect 5724 2586 5776 2592
rect 6656 2514 6684 2604
rect 6828 2586 6880 2592
rect 6644 2508 6696 2514
rect 6644 2450 6696 2456
rect 7208 2446 7236 2746
rect 8036 2650 8064 2926
rect 8114 2748 8422 2757
rect 8114 2746 8120 2748
rect 8176 2746 8200 2748
rect 8256 2746 8280 2748
rect 8336 2746 8360 2748
rect 8416 2746 8422 2748
rect 8176 2694 8178 2746
rect 8358 2694 8360 2746
rect 8114 2692 8120 2694
rect 8176 2692 8200 2694
rect 8256 2692 8280 2694
rect 8336 2692 8360 2694
rect 8416 2692 8422 2694
rect 8114 2683 8422 2692
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 5172 2372 5224 2378
rect 5172 2314 5224 2320
rect 2504 2304 2556 2310
rect 2504 2246 2556 2252
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 2633 2204 2941 2213
rect 2633 2202 2639 2204
rect 2695 2202 2719 2204
rect 2775 2202 2799 2204
rect 2855 2202 2879 2204
rect 2935 2202 2941 2204
rect 2695 2150 2697 2202
rect 2877 2150 2879 2202
rect 2633 2148 2639 2150
rect 2695 2148 2719 2150
rect 2775 2148 2799 2150
rect 2855 2148 2879 2150
rect 2935 2148 2941 2150
rect 2633 2139 2941 2148
rect 4680 2204 4988 2213
rect 4680 2202 4686 2204
rect 4742 2202 4766 2204
rect 4822 2202 4846 2204
rect 4902 2202 4926 2204
rect 4982 2202 4988 2204
rect 4742 2150 4744 2202
rect 4924 2150 4926 2202
rect 4680 2148 4686 2150
rect 4742 2148 4766 2150
rect 4822 2148 4846 2150
rect 4902 2148 4926 2150
rect 4982 2148 4988 2150
rect 4680 2139 4988 2148
rect 5184 800 5212 2314
rect 6727 2204 7035 2213
rect 6727 2202 6733 2204
rect 6789 2202 6813 2204
rect 6869 2202 6893 2204
rect 6949 2202 6973 2204
rect 7029 2202 7035 2204
rect 6789 2150 6791 2202
rect 6971 2150 6973 2202
rect 6727 2148 6733 2150
rect 6789 2148 6813 2150
rect 6869 2148 6893 2150
rect 6949 2148 6973 2150
rect 7029 2148 7035 2150
rect 6727 2139 7035 2148
rect 8774 2204 9082 2213
rect 8774 2202 8780 2204
rect 8836 2202 8860 2204
rect 8916 2202 8940 2204
rect 8996 2202 9020 2204
rect 9076 2202 9082 2204
rect 8836 2150 8838 2202
rect 9018 2150 9020 2202
rect 8774 2148 8780 2150
rect 8836 2148 8860 2150
rect 8916 2148 8940 2150
rect 8996 2148 9020 2150
rect 9076 2148 9082 2150
rect 8774 2139 9082 2148
rect 5170 0 5226 800
<< via2 >>
rect 1979 10362 2035 10364
rect 2059 10362 2115 10364
rect 2139 10362 2195 10364
rect 2219 10362 2275 10364
rect 1979 10310 2025 10362
rect 2025 10310 2035 10362
rect 2059 10310 2089 10362
rect 2089 10310 2101 10362
rect 2101 10310 2115 10362
rect 2139 10310 2153 10362
rect 2153 10310 2165 10362
rect 2165 10310 2195 10362
rect 2219 10310 2229 10362
rect 2229 10310 2275 10362
rect 1979 10308 2035 10310
rect 2059 10308 2115 10310
rect 2139 10308 2195 10310
rect 2219 10308 2275 10310
rect 4026 10362 4082 10364
rect 4106 10362 4162 10364
rect 4186 10362 4242 10364
rect 4266 10362 4322 10364
rect 4026 10310 4072 10362
rect 4072 10310 4082 10362
rect 4106 10310 4136 10362
rect 4136 10310 4148 10362
rect 4148 10310 4162 10362
rect 4186 10310 4200 10362
rect 4200 10310 4212 10362
rect 4212 10310 4242 10362
rect 4266 10310 4276 10362
rect 4276 10310 4322 10362
rect 4026 10308 4082 10310
rect 4106 10308 4162 10310
rect 4186 10308 4242 10310
rect 4266 10308 4322 10310
rect 6073 10362 6129 10364
rect 6153 10362 6209 10364
rect 6233 10362 6289 10364
rect 6313 10362 6369 10364
rect 6073 10310 6119 10362
rect 6119 10310 6129 10362
rect 6153 10310 6183 10362
rect 6183 10310 6195 10362
rect 6195 10310 6209 10362
rect 6233 10310 6247 10362
rect 6247 10310 6259 10362
rect 6259 10310 6289 10362
rect 6313 10310 6323 10362
rect 6323 10310 6369 10362
rect 6073 10308 6129 10310
rect 6153 10308 6209 10310
rect 6233 10308 6289 10310
rect 6313 10308 6369 10310
rect 8120 10362 8176 10364
rect 8200 10362 8256 10364
rect 8280 10362 8336 10364
rect 8360 10362 8416 10364
rect 8120 10310 8166 10362
rect 8166 10310 8176 10362
rect 8200 10310 8230 10362
rect 8230 10310 8242 10362
rect 8242 10310 8256 10362
rect 8280 10310 8294 10362
rect 8294 10310 8306 10362
rect 8306 10310 8336 10362
rect 8360 10310 8370 10362
rect 8370 10310 8416 10362
rect 8120 10308 8176 10310
rect 8200 10308 8256 10310
rect 8280 10308 8336 10310
rect 8360 10308 8416 10310
rect 1582 8880 1638 8936
rect 1306 6160 1362 6216
rect 1979 9274 2035 9276
rect 2059 9274 2115 9276
rect 2139 9274 2195 9276
rect 2219 9274 2275 9276
rect 1979 9222 2025 9274
rect 2025 9222 2035 9274
rect 2059 9222 2089 9274
rect 2089 9222 2101 9274
rect 2101 9222 2115 9274
rect 2139 9222 2153 9274
rect 2153 9222 2165 9274
rect 2165 9222 2195 9274
rect 2219 9222 2229 9274
rect 2229 9222 2275 9274
rect 1979 9220 2035 9222
rect 2059 9220 2115 9222
rect 2139 9220 2195 9222
rect 2219 9220 2275 9222
rect 1858 8356 1914 8392
rect 1858 8336 1860 8356
rect 1860 8336 1912 8356
rect 1912 8336 1914 8356
rect 2639 9818 2695 9820
rect 2719 9818 2775 9820
rect 2799 9818 2855 9820
rect 2879 9818 2935 9820
rect 2639 9766 2685 9818
rect 2685 9766 2695 9818
rect 2719 9766 2749 9818
rect 2749 9766 2761 9818
rect 2761 9766 2775 9818
rect 2799 9766 2813 9818
rect 2813 9766 2825 9818
rect 2825 9766 2855 9818
rect 2879 9766 2889 9818
rect 2889 9766 2935 9818
rect 2639 9764 2695 9766
rect 2719 9764 2775 9766
rect 2799 9764 2855 9766
rect 2879 9764 2935 9766
rect 2639 8730 2695 8732
rect 2719 8730 2775 8732
rect 2799 8730 2855 8732
rect 2879 8730 2935 8732
rect 2639 8678 2685 8730
rect 2685 8678 2695 8730
rect 2719 8678 2749 8730
rect 2749 8678 2761 8730
rect 2761 8678 2775 8730
rect 2799 8678 2813 8730
rect 2813 8678 2825 8730
rect 2825 8678 2855 8730
rect 2879 8678 2889 8730
rect 2889 8678 2935 8730
rect 2639 8676 2695 8678
rect 2719 8676 2775 8678
rect 2799 8676 2855 8678
rect 2879 8676 2935 8678
rect 1979 8186 2035 8188
rect 2059 8186 2115 8188
rect 2139 8186 2195 8188
rect 2219 8186 2275 8188
rect 1979 8134 2025 8186
rect 2025 8134 2035 8186
rect 2059 8134 2089 8186
rect 2089 8134 2101 8186
rect 2101 8134 2115 8186
rect 2139 8134 2153 8186
rect 2153 8134 2165 8186
rect 2165 8134 2195 8186
rect 2219 8134 2229 8186
rect 2229 8134 2275 8186
rect 1979 8132 2035 8134
rect 2059 8132 2115 8134
rect 2139 8132 2195 8134
rect 2219 8132 2275 8134
rect 2318 7812 2374 7848
rect 2318 7792 2320 7812
rect 2320 7792 2372 7812
rect 2372 7792 2374 7812
rect 1979 7098 2035 7100
rect 2059 7098 2115 7100
rect 2139 7098 2195 7100
rect 2219 7098 2275 7100
rect 1979 7046 2025 7098
rect 2025 7046 2035 7098
rect 2059 7046 2089 7098
rect 2089 7046 2101 7098
rect 2101 7046 2115 7098
rect 2139 7046 2153 7098
rect 2153 7046 2165 7098
rect 2165 7046 2195 7098
rect 2219 7046 2229 7098
rect 2229 7046 2275 7098
rect 1979 7044 2035 7046
rect 2059 7044 2115 7046
rect 2139 7044 2195 7046
rect 2219 7044 2275 7046
rect 2962 7928 3018 7984
rect 2639 7642 2695 7644
rect 2719 7642 2775 7644
rect 2799 7642 2855 7644
rect 2879 7642 2935 7644
rect 2639 7590 2685 7642
rect 2685 7590 2695 7642
rect 2719 7590 2749 7642
rect 2749 7590 2761 7642
rect 2761 7590 2775 7642
rect 2799 7590 2813 7642
rect 2813 7590 2825 7642
rect 2825 7590 2855 7642
rect 2879 7590 2889 7642
rect 2889 7590 2935 7642
rect 2639 7588 2695 7590
rect 2719 7588 2775 7590
rect 2799 7588 2855 7590
rect 2879 7588 2935 7590
rect 1950 6840 2006 6896
rect 2639 6554 2695 6556
rect 2719 6554 2775 6556
rect 2799 6554 2855 6556
rect 2879 6554 2935 6556
rect 2639 6502 2685 6554
rect 2685 6502 2695 6554
rect 2719 6502 2749 6554
rect 2749 6502 2761 6554
rect 2761 6502 2775 6554
rect 2799 6502 2813 6554
rect 2813 6502 2825 6554
rect 2825 6502 2855 6554
rect 2879 6502 2889 6554
rect 2889 6502 2935 6554
rect 2639 6500 2695 6502
rect 2719 6500 2775 6502
rect 2799 6500 2855 6502
rect 2879 6500 2935 6502
rect 1582 6160 1638 6216
rect 1979 6010 2035 6012
rect 2059 6010 2115 6012
rect 2139 6010 2195 6012
rect 2219 6010 2275 6012
rect 1979 5958 2025 6010
rect 2025 5958 2035 6010
rect 2059 5958 2089 6010
rect 2089 5958 2101 6010
rect 2101 5958 2115 6010
rect 2139 5958 2153 6010
rect 2153 5958 2165 6010
rect 2165 5958 2195 6010
rect 2219 5958 2229 6010
rect 2229 5958 2275 6010
rect 1979 5956 2035 5958
rect 2059 5956 2115 5958
rect 2139 5956 2195 5958
rect 2219 5956 2275 5958
rect 1766 5208 1822 5264
rect 1979 4922 2035 4924
rect 2059 4922 2115 4924
rect 2139 4922 2195 4924
rect 2219 4922 2275 4924
rect 1979 4870 2025 4922
rect 2025 4870 2035 4922
rect 2059 4870 2089 4922
rect 2089 4870 2101 4922
rect 2101 4870 2115 4922
rect 2139 4870 2153 4922
rect 2153 4870 2165 4922
rect 2165 4870 2195 4922
rect 2219 4870 2229 4922
rect 2229 4870 2275 4922
rect 1979 4868 2035 4870
rect 2059 4868 2115 4870
rect 2139 4868 2195 4870
rect 2219 4868 2275 4870
rect 2870 5616 2926 5672
rect 2639 5466 2695 5468
rect 2719 5466 2775 5468
rect 2799 5466 2855 5468
rect 2879 5466 2935 5468
rect 2639 5414 2685 5466
rect 2685 5414 2695 5466
rect 2719 5414 2749 5466
rect 2749 5414 2761 5466
rect 2761 5414 2775 5466
rect 2799 5414 2813 5466
rect 2813 5414 2825 5466
rect 2825 5414 2855 5466
rect 2879 5414 2889 5466
rect 2889 5414 2935 5466
rect 2639 5412 2695 5414
rect 2719 5412 2775 5414
rect 2799 5412 2855 5414
rect 2879 5412 2935 5414
rect 4434 9560 4490 9616
rect 4686 9818 4742 9820
rect 4766 9818 4822 9820
rect 4846 9818 4902 9820
rect 4926 9818 4982 9820
rect 4686 9766 4732 9818
rect 4732 9766 4742 9818
rect 4766 9766 4796 9818
rect 4796 9766 4808 9818
rect 4808 9766 4822 9818
rect 4846 9766 4860 9818
rect 4860 9766 4872 9818
rect 4872 9766 4902 9818
rect 4926 9766 4936 9818
rect 4936 9766 4982 9818
rect 4686 9764 4742 9766
rect 4766 9764 4822 9766
rect 4846 9764 4902 9766
rect 4926 9764 4982 9766
rect 4026 9274 4082 9276
rect 4106 9274 4162 9276
rect 4186 9274 4242 9276
rect 4266 9274 4322 9276
rect 4026 9222 4072 9274
rect 4072 9222 4082 9274
rect 4106 9222 4136 9274
rect 4136 9222 4148 9274
rect 4148 9222 4162 9274
rect 4186 9222 4200 9274
rect 4200 9222 4212 9274
rect 4212 9222 4242 9274
rect 4266 9222 4276 9274
rect 4276 9222 4322 9274
rect 4026 9220 4082 9222
rect 4106 9220 4162 9222
rect 4186 9220 4242 9222
rect 4266 9220 4322 9222
rect 3974 8880 4030 8936
rect 3330 7928 3386 7984
rect 3606 8336 3662 8392
rect 3606 7828 3608 7848
rect 3608 7828 3660 7848
rect 3660 7828 3662 7848
rect 3606 7792 3662 7828
rect 3238 6568 3294 6624
rect 3238 6432 3294 6488
rect 3514 6704 3570 6760
rect 1979 3834 2035 3836
rect 2059 3834 2115 3836
rect 2139 3834 2195 3836
rect 2219 3834 2275 3836
rect 1979 3782 2025 3834
rect 2025 3782 2035 3834
rect 2059 3782 2089 3834
rect 2089 3782 2101 3834
rect 2101 3782 2115 3834
rect 2139 3782 2153 3834
rect 2153 3782 2165 3834
rect 2165 3782 2195 3834
rect 2219 3782 2229 3834
rect 2229 3782 2275 3834
rect 1979 3780 2035 3782
rect 2059 3780 2115 3782
rect 2139 3780 2195 3782
rect 2219 3780 2275 3782
rect 2410 3984 2466 4040
rect 2639 4378 2695 4380
rect 2719 4378 2775 4380
rect 2799 4378 2855 4380
rect 2879 4378 2935 4380
rect 2639 4326 2685 4378
rect 2685 4326 2695 4378
rect 2719 4326 2749 4378
rect 2749 4326 2761 4378
rect 2761 4326 2775 4378
rect 2799 4326 2813 4378
rect 2813 4326 2825 4378
rect 2825 4326 2855 4378
rect 2879 4326 2889 4378
rect 2889 4326 2935 4378
rect 2639 4324 2695 4326
rect 2719 4324 2775 4326
rect 2799 4324 2855 4326
rect 2879 4324 2935 4326
rect 3330 5616 3386 5672
rect 1979 2746 2035 2748
rect 2059 2746 2115 2748
rect 2139 2746 2195 2748
rect 2219 2746 2275 2748
rect 1979 2694 2025 2746
rect 2025 2694 2035 2746
rect 2059 2694 2089 2746
rect 2089 2694 2101 2746
rect 2101 2694 2115 2746
rect 2139 2694 2153 2746
rect 2153 2694 2165 2746
rect 2165 2694 2195 2746
rect 2219 2694 2229 2746
rect 2229 2694 2275 2746
rect 1979 2692 2035 2694
rect 2059 2692 2115 2694
rect 2139 2692 2195 2694
rect 2219 2692 2275 2694
rect 2639 3290 2695 3292
rect 2719 3290 2775 3292
rect 2799 3290 2855 3292
rect 2879 3290 2935 3292
rect 2639 3238 2685 3290
rect 2685 3238 2695 3290
rect 2719 3238 2749 3290
rect 2749 3238 2761 3290
rect 2761 3238 2775 3290
rect 2799 3238 2813 3290
rect 2813 3238 2825 3290
rect 2825 3238 2855 3290
rect 2879 3238 2889 3290
rect 2889 3238 2935 3290
rect 2639 3236 2695 3238
rect 2719 3236 2775 3238
rect 2799 3236 2855 3238
rect 2879 3236 2935 3238
rect 4026 8186 4082 8188
rect 4106 8186 4162 8188
rect 4186 8186 4242 8188
rect 4266 8186 4322 8188
rect 4026 8134 4072 8186
rect 4072 8134 4082 8186
rect 4106 8134 4136 8186
rect 4136 8134 4148 8186
rect 4148 8134 4162 8186
rect 4186 8134 4200 8186
rect 4200 8134 4212 8186
rect 4212 8134 4242 8186
rect 4266 8134 4276 8186
rect 4276 8134 4322 8186
rect 4026 8132 4082 8134
rect 4106 8132 4162 8134
rect 4186 8132 4242 8134
rect 4266 8132 4322 8134
rect 4026 7098 4082 7100
rect 4106 7098 4162 7100
rect 4186 7098 4242 7100
rect 4266 7098 4322 7100
rect 4026 7046 4072 7098
rect 4072 7046 4082 7098
rect 4106 7046 4136 7098
rect 4136 7046 4148 7098
rect 4148 7046 4162 7098
rect 4186 7046 4200 7098
rect 4200 7046 4212 7098
rect 4212 7046 4242 7098
rect 4266 7046 4276 7098
rect 4276 7046 4322 7098
rect 4026 7044 4082 7046
rect 4106 7044 4162 7046
rect 4186 7044 4242 7046
rect 4266 7044 4322 7046
rect 3790 6704 3846 6760
rect 3698 6568 3754 6624
rect 4066 6704 4122 6760
rect 3974 6432 4030 6488
rect 3974 6196 3976 6216
rect 3976 6196 4028 6216
rect 4028 6196 4030 6216
rect 3974 6160 4030 6196
rect 4686 8730 4742 8732
rect 4766 8730 4822 8732
rect 4846 8730 4902 8732
rect 4926 8730 4982 8732
rect 4686 8678 4732 8730
rect 4732 8678 4742 8730
rect 4766 8678 4796 8730
rect 4796 8678 4808 8730
rect 4808 8678 4822 8730
rect 4846 8678 4860 8730
rect 4860 8678 4872 8730
rect 4872 8678 4902 8730
rect 4926 8678 4936 8730
rect 4936 8678 4982 8730
rect 4686 8676 4742 8678
rect 4766 8676 4822 8678
rect 4846 8676 4902 8678
rect 4926 8676 4982 8678
rect 4686 7642 4742 7644
rect 4766 7642 4822 7644
rect 4846 7642 4902 7644
rect 4926 7642 4982 7644
rect 4686 7590 4732 7642
rect 4732 7590 4742 7642
rect 4766 7590 4796 7642
rect 4796 7590 4808 7642
rect 4808 7590 4822 7642
rect 4846 7590 4860 7642
rect 4860 7590 4872 7642
rect 4872 7590 4902 7642
rect 4926 7590 4936 7642
rect 4936 7590 4982 7642
rect 4686 7588 4742 7590
rect 4766 7588 4822 7590
rect 4846 7588 4902 7590
rect 4926 7588 4982 7590
rect 4986 7384 5042 7440
rect 4986 6976 5042 7032
rect 4894 6840 4950 6896
rect 4026 6010 4082 6012
rect 4106 6010 4162 6012
rect 4186 6010 4242 6012
rect 4266 6010 4322 6012
rect 4026 5958 4072 6010
rect 4072 5958 4082 6010
rect 4106 5958 4136 6010
rect 4136 5958 4148 6010
rect 4148 5958 4162 6010
rect 4186 5958 4200 6010
rect 4200 5958 4212 6010
rect 4212 5958 4242 6010
rect 4266 5958 4276 6010
rect 4276 5958 4322 6010
rect 4026 5956 4082 5958
rect 4106 5956 4162 5958
rect 4186 5956 4242 5958
rect 4266 5956 4322 5958
rect 4026 4922 4082 4924
rect 4106 4922 4162 4924
rect 4186 4922 4242 4924
rect 4266 4922 4322 4924
rect 4026 4870 4072 4922
rect 4072 4870 4082 4922
rect 4106 4870 4136 4922
rect 4136 4870 4148 4922
rect 4148 4870 4162 4922
rect 4186 4870 4200 4922
rect 4200 4870 4212 4922
rect 4212 4870 4242 4922
rect 4266 4870 4276 4922
rect 4276 4870 4322 4922
rect 4026 4868 4082 4870
rect 4106 4868 4162 4870
rect 4186 4868 4242 4870
rect 4266 4868 4322 4870
rect 4686 6554 4742 6556
rect 4766 6554 4822 6556
rect 4846 6554 4902 6556
rect 4926 6554 4982 6556
rect 4686 6502 4732 6554
rect 4732 6502 4742 6554
rect 4766 6502 4796 6554
rect 4796 6502 4808 6554
rect 4808 6502 4822 6554
rect 4846 6502 4860 6554
rect 4860 6502 4872 6554
rect 4872 6502 4902 6554
rect 4926 6502 4936 6554
rect 4936 6502 4982 6554
rect 4686 6500 4742 6502
rect 4766 6500 4822 6502
rect 4846 6500 4902 6502
rect 4926 6500 4982 6502
rect 4686 5466 4742 5468
rect 4766 5466 4822 5468
rect 4846 5466 4902 5468
rect 4926 5466 4982 5468
rect 4686 5414 4732 5466
rect 4732 5414 4742 5466
rect 4766 5414 4796 5466
rect 4796 5414 4808 5466
rect 4808 5414 4822 5466
rect 4846 5414 4860 5466
rect 4860 5414 4872 5466
rect 4872 5414 4902 5466
rect 4926 5414 4936 5466
rect 4936 5414 4982 5466
rect 4686 5412 4742 5414
rect 4766 5412 4822 5414
rect 4846 5412 4902 5414
rect 4926 5412 4982 5414
rect 6733 9818 6789 9820
rect 6813 9818 6869 9820
rect 6893 9818 6949 9820
rect 6973 9818 7029 9820
rect 6733 9766 6779 9818
rect 6779 9766 6789 9818
rect 6813 9766 6843 9818
rect 6843 9766 6855 9818
rect 6855 9766 6869 9818
rect 6893 9766 6907 9818
rect 6907 9766 6919 9818
rect 6919 9766 6949 9818
rect 6973 9766 6983 9818
rect 6983 9766 7029 9818
rect 6733 9764 6789 9766
rect 6813 9764 6869 9766
rect 6893 9764 6949 9766
rect 6973 9764 7029 9766
rect 6073 9274 6129 9276
rect 6153 9274 6209 9276
rect 6233 9274 6289 9276
rect 6313 9274 6369 9276
rect 6073 9222 6119 9274
rect 6119 9222 6129 9274
rect 6153 9222 6183 9274
rect 6183 9222 6195 9274
rect 6195 9222 6209 9274
rect 6233 9222 6247 9274
rect 6247 9222 6259 9274
rect 6259 9222 6289 9274
rect 6313 9222 6323 9274
rect 6323 9222 6369 9274
rect 6073 9220 6129 9222
rect 6153 9220 6209 9222
rect 6233 9220 6289 9222
rect 6313 9220 6369 9222
rect 5354 7540 5410 7576
rect 5354 7520 5356 7540
rect 5356 7520 5408 7540
rect 5408 7520 5410 7540
rect 6182 8916 6184 8936
rect 6184 8916 6236 8936
rect 6236 8916 6238 8936
rect 6182 8880 6238 8916
rect 6073 8186 6129 8188
rect 6153 8186 6209 8188
rect 6233 8186 6289 8188
rect 6313 8186 6369 8188
rect 6073 8134 6119 8186
rect 6119 8134 6129 8186
rect 6153 8134 6183 8186
rect 6183 8134 6195 8186
rect 6195 8134 6209 8186
rect 6233 8134 6247 8186
rect 6247 8134 6259 8186
rect 6259 8134 6289 8186
rect 6313 8134 6323 8186
rect 6323 8134 6369 8186
rect 6073 8132 6129 8134
rect 6153 8132 6209 8134
rect 6233 8132 6289 8134
rect 6313 8132 6369 8134
rect 5354 5652 5356 5672
rect 5356 5652 5408 5672
rect 5408 5652 5410 5672
rect 5354 5616 5410 5652
rect 4434 4564 4436 4584
rect 4436 4564 4488 4584
rect 4488 4564 4490 4584
rect 4434 4528 4490 4564
rect 4026 3834 4082 3836
rect 4106 3834 4162 3836
rect 4186 3834 4242 3836
rect 4266 3834 4322 3836
rect 4026 3782 4072 3834
rect 4072 3782 4082 3834
rect 4106 3782 4136 3834
rect 4136 3782 4148 3834
rect 4148 3782 4162 3834
rect 4186 3782 4200 3834
rect 4200 3782 4212 3834
rect 4212 3782 4242 3834
rect 4266 3782 4276 3834
rect 4276 3782 4322 3834
rect 4026 3780 4082 3782
rect 4106 3780 4162 3782
rect 4186 3780 4242 3782
rect 4266 3780 4322 3782
rect 4686 4378 4742 4380
rect 4766 4378 4822 4380
rect 4846 4378 4902 4380
rect 4926 4378 4982 4380
rect 4686 4326 4732 4378
rect 4732 4326 4742 4378
rect 4766 4326 4796 4378
rect 4796 4326 4808 4378
rect 4808 4326 4822 4378
rect 4846 4326 4860 4378
rect 4860 4326 4872 4378
rect 4872 4326 4902 4378
rect 4926 4326 4936 4378
rect 4936 4326 4982 4378
rect 4686 4324 4742 4326
rect 4766 4324 4822 4326
rect 4846 4324 4902 4326
rect 4926 4324 4982 4326
rect 4026 2746 4082 2748
rect 4106 2746 4162 2748
rect 4186 2746 4242 2748
rect 4266 2746 4322 2748
rect 4026 2694 4072 2746
rect 4072 2694 4082 2746
rect 4106 2694 4136 2746
rect 4136 2694 4148 2746
rect 4148 2694 4162 2746
rect 4186 2694 4200 2746
rect 4200 2694 4212 2746
rect 4212 2694 4242 2746
rect 4266 2694 4276 2746
rect 4276 2694 4322 2746
rect 4026 2692 4082 2694
rect 4106 2692 4162 2694
rect 4186 2692 4242 2694
rect 4266 2692 4322 2694
rect 4710 3476 4712 3496
rect 4712 3476 4764 3496
rect 4764 3476 4766 3496
rect 4710 3440 4766 3476
rect 5998 7384 6054 7440
rect 6733 8730 6789 8732
rect 6813 8730 6869 8732
rect 6893 8730 6949 8732
rect 6973 8730 7029 8732
rect 6733 8678 6779 8730
rect 6779 8678 6789 8730
rect 6813 8678 6843 8730
rect 6843 8678 6855 8730
rect 6855 8678 6869 8730
rect 6893 8678 6907 8730
rect 6907 8678 6919 8730
rect 6919 8678 6949 8730
rect 6973 8678 6983 8730
rect 6983 8678 7029 8730
rect 6733 8676 6789 8678
rect 6813 8676 6869 8678
rect 6893 8676 6949 8678
rect 6973 8676 7029 8678
rect 8780 9818 8836 9820
rect 8860 9818 8916 9820
rect 8940 9818 8996 9820
rect 9020 9818 9076 9820
rect 8780 9766 8826 9818
rect 8826 9766 8836 9818
rect 8860 9766 8890 9818
rect 8890 9766 8902 9818
rect 8902 9766 8916 9818
rect 8940 9766 8954 9818
rect 8954 9766 8966 9818
rect 8966 9766 8996 9818
rect 9020 9766 9030 9818
rect 9030 9766 9076 9818
rect 8780 9764 8836 9766
rect 8860 9764 8916 9766
rect 8940 9764 8996 9766
rect 9020 9764 9076 9766
rect 7562 8880 7618 8936
rect 6733 7642 6789 7644
rect 6813 7642 6869 7644
rect 6893 7642 6949 7644
rect 6973 7642 7029 7644
rect 6733 7590 6779 7642
rect 6779 7590 6789 7642
rect 6813 7590 6843 7642
rect 6843 7590 6855 7642
rect 6855 7590 6869 7642
rect 6893 7590 6907 7642
rect 6907 7590 6919 7642
rect 6919 7590 6949 7642
rect 6973 7590 6983 7642
rect 6983 7590 7029 7642
rect 6733 7588 6789 7590
rect 6813 7588 6869 7590
rect 6893 7588 6949 7590
rect 6973 7588 7029 7590
rect 6073 7098 6129 7100
rect 6153 7098 6209 7100
rect 6233 7098 6289 7100
rect 6313 7098 6369 7100
rect 6073 7046 6119 7098
rect 6119 7046 6129 7098
rect 6153 7046 6183 7098
rect 6183 7046 6195 7098
rect 6195 7046 6209 7098
rect 6233 7046 6247 7098
rect 6247 7046 6259 7098
rect 6259 7046 6289 7098
rect 6313 7046 6323 7098
rect 6323 7046 6369 7098
rect 6073 7044 6129 7046
rect 6153 7044 6209 7046
rect 6233 7044 6289 7046
rect 6313 7044 6369 7046
rect 6182 6840 6238 6896
rect 6366 6160 6422 6216
rect 6826 6740 6828 6760
rect 6828 6740 6880 6760
rect 6880 6740 6882 6760
rect 6826 6704 6882 6740
rect 6733 6554 6789 6556
rect 6813 6554 6869 6556
rect 6893 6554 6949 6556
rect 6973 6554 7029 6556
rect 6733 6502 6779 6554
rect 6779 6502 6789 6554
rect 6813 6502 6843 6554
rect 6843 6502 6855 6554
rect 6855 6502 6869 6554
rect 6893 6502 6907 6554
rect 6907 6502 6919 6554
rect 6919 6502 6949 6554
rect 6973 6502 6983 6554
rect 6983 6502 7029 6554
rect 6733 6500 6789 6502
rect 6813 6500 6869 6502
rect 6893 6500 6949 6502
rect 6973 6500 7029 6502
rect 6073 6010 6129 6012
rect 6153 6010 6209 6012
rect 6233 6010 6289 6012
rect 6313 6010 6369 6012
rect 6073 5958 6119 6010
rect 6119 5958 6129 6010
rect 6153 5958 6183 6010
rect 6183 5958 6195 6010
rect 6195 5958 6209 6010
rect 6233 5958 6247 6010
rect 6247 5958 6259 6010
rect 6259 5958 6289 6010
rect 6313 5958 6323 6010
rect 6323 5958 6369 6010
rect 6073 5956 6129 5958
rect 6153 5956 6209 5958
rect 6233 5956 6289 5958
rect 6313 5956 6369 5958
rect 5722 4564 5724 4584
rect 5724 4564 5776 4584
rect 5776 4564 5778 4584
rect 5722 4528 5778 4564
rect 6274 5208 6330 5264
rect 6734 6160 6790 6216
rect 7286 7404 7342 7440
rect 7286 7384 7288 7404
rect 7288 7384 7340 7404
rect 7340 7384 7342 7404
rect 8120 9274 8176 9276
rect 8200 9274 8256 9276
rect 8280 9274 8336 9276
rect 8360 9274 8416 9276
rect 8120 9222 8166 9274
rect 8166 9222 8176 9274
rect 8200 9222 8230 9274
rect 8230 9222 8242 9274
rect 8242 9222 8256 9274
rect 8280 9222 8294 9274
rect 8294 9222 8306 9274
rect 8306 9222 8336 9274
rect 8360 9222 8370 9274
rect 8370 9222 8416 9274
rect 8120 9220 8176 9222
rect 8200 9220 8256 9222
rect 8280 9220 8336 9222
rect 8360 9220 8416 9222
rect 8780 8730 8836 8732
rect 8860 8730 8916 8732
rect 8940 8730 8996 8732
rect 9020 8730 9076 8732
rect 8780 8678 8826 8730
rect 8826 8678 8836 8730
rect 8860 8678 8890 8730
rect 8890 8678 8902 8730
rect 8902 8678 8916 8730
rect 8940 8678 8954 8730
rect 8954 8678 8966 8730
rect 8966 8678 8996 8730
rect 9020 8678 9030 8730
rect 9030 8678 9076 8730
rect 8780 8676 8836 8678
rect 8860 8676 8916 8678
rect 8940 8676 8996 8678
rect 9020 8676 9076 8678
rect 8120 8186 8176 8188
rect 8200 8186 8256 8188
rect 8280 8186 8336 8188
rect 8360 8186 8416 8188
rect 8120 8134 8166 8186
rect 8166 8134 8176 8186
rect 8200 8134 8230 8186
rect 8230 8134 8242 8186
rect 8242 8134 8256 8186
rect 8280 8134 8294 8186
rect 8294 8134 8306 8186
rect 8306 8134 8336 8186
rect 8360 8134 8370 8186
rect 8370 8134 8416 8186
rect 8120 8132 8176 8134
rect 8200 8132 8256 8134
rect 8280 8132 8336 8134
rect 8360 8132 8416 8134
rect 6733 5466 6789 5468
rect 6813 5466 6869 5468
rect 6893 5466 6949 5468
rect 6973 5466 7029 5468
rect 6733 5414 6779 5466
rect 6779 5414 6789 5466
rect 6813 5414 6843 5466
rect 6843 5414 6855 5466
rect 6855 5414 6869 5466
rect 6893 5414 6907 5466
rect 6907 5414 6919 5466
rect 6919 5414 6949 5466
rect 6973 5414 6983 5466
rect 6983 5414 7029 5466
rect 6733 5412 6789 5414
rect 6813 5412 6869 5414
rect 6893 5412 6949 5414
rect 6973 5412 7029 5414
rect 6073 4922 6129 4924
rect 6153 4922 6209 4924
rect 6233 4922 6289 4924
rect 6313 4922 6369 4924
rect 6073 4870 6119 4922
rect 6119 4870 6129 4922
rect 6153 4870 6183 4922
rect 6183 4870 6195 4922
rect 6195 4870 6209 4922
rect 6233 4870 6247 4922
rect 6247 4870 6259 4922
rect 6259 4870 6289 4922
rect 6313 4870 6323 4922
rect 6323 4870 6369 4922
rect 6073 4868 6129 4870
rect 6153 4868 6209 4870
rect 6233 4868 6289 4870
rect 6313 4868 6369 4870
rect 6274 4664 6330 4720
rect 5630 3984 5686 4040
rect 5538 3476 5540 3496
rect 5540 3476 5592 3496
rect 5592 3476 5594 3496
rect 4686 3290 4742 3292
rect 4766 3290 4822 3292
rect 4846 3290 4902 3292
rect 4926 3290 4982 3292
rect 4686 3238 4732 3290
rect 4732 3238 4742 3290
rect 4766 3238 4796 3290
rect 4796 3238 4808 3290
rect 4808 3238 4822 3290
rect 4846 3238 4860 3290
rect 4860 3238 4872 3290
rect 4872 3238 4902 3290
rect 4926 3238 4936 3290
rect 4936 3238 4982 3290
rect 4686 3236 4742 3238
rect 4766 3236 4822 3238
rect 4846 3236 4902 3238
rect 4926 3236 4982 3238
rect 5538 3440 5594 3476
rect 6073 3834 6129 3836
rect 6153 3834 6209 3836
rect 6233 3834 6289 3836
rect 6313 3834 6369 3836
rect 6073 3782 6119 3834
rect 6119 3782 6129 3834
rect 6153 3782 6183 3834
rect 6183 3782 6195 3834
rect 6195 3782 6209 3834
rect 6233 3782 6247 3834
rect 6247 3782 6259 3834
rect 6259 3782 6289 3834
rect 6313 3782 6323 3834
rect 6323 3782 6369 3834
rect 6073 3780 6129 3782
rect 6153 3780 6209 3782
rect 6233 3780 6289 3782
rect 6313 3780 6369 3782
rect 6073 2746 6129 2748
rect 6153 2746 6209 2748
rect 6233 2746 6289 2748
rect 6313 2746 6369 2748
rect 6073 2694 6119 2746
rect 6119 2694 6129 2746
rect 6153 2694 6183 2746
rect 6183 2694 6195 2746
rect 6195 2694 6209 2746
rect 6233 2694 6247 2746
rect 6247 2694 6259 2746
rect 6259 2694 6289 2746
rect 6313 2694 6323 2746
rect 6323 2694 6369 2746
rect 6073 2692 6129 2694
rect 6153 2692 6209 2694
rect 6233 2692 6289 2694
rect 6313 2692 6369 2694
rect 7470 5616 7526 5672
rect 8780 7642 8836 7644
rect 8860 7642 8916 7644
rect 8940 7642 8996 7644
rect 9020 7642 9076 7644
rect 8780 7590 8826 7642
rect 8826 7590 8836 7642
rect 8860 7590 8890 7642
rect 8890 7590 8902 7642
rect 8902 7590 8916 7642
rect 8940 7590 8954 7642
rect 8954 7590 8966 7642
rect 8966 7590 8996 7642
rect 9020 7590 9030 7642
rect 9030 7590 9076 7642
rect 8780 7588 8836 7590
rect 8860 7588 8916 7590
rect 8940 7588 8996 7590
rect 9020 7588 9076 7590
rect 8120 7098 8176 7100
rect 8200 7098 8256 7100
rect 8280 7098 8336 7100
rect 8360 7098 8416 7100
rect 8120 7046 8166 7098
rect 8166 7046 8176 7098
rect 8200 7046 8230 7098
rect 8230 7046 8242 7098
rect 8242 7046 8256 7098
rect 8280 7046 8294 7098
rect 8294 7046 8306 7098
rect 8306 7046 8336 7098
rect 8360 7046 8370 7098
rect 8370 7046 8416 7098
rect 8120 7044 8176 7046
rect 8200 7044 8256 7046
rect 8280 7044 8336 7046
rect 8360 7044 8416 7046
rect 8120 6010 8176 6012
rect 8200 6010 8256 6012
rect 8280 6010 8336 6012
rect 8360 6010 8416 6012
rect 8120 5958 8166 6010
rect 8166 5958 8176 6010
rect 8200 5958 8230 6010
rect 8230 5958 8242 6010
rect 8242 5958 8256 6010
rect 8280 5958 8294 6010
rect 8294 5958 8306 6010
rect 8306 5958 8336 6010
rect 8360 5958 8370 6010
rect 8370 5958 8416 6010
rect 8120 5956 8176 5958
rect 8200 5956 8256 5958
rect 8280 5956 8336 5958
rect 8360 5956 8416 5958
rect 6733 4378 6789 4380
rect 6813 4378 6869 4380
rect 6893 4378 6949 4380
rect 6973 4378 7029 4380
rect 6733 4326 6779 4378
rect 6779 4326 6789 4378
rect 6813 4326 6843 4378
rect 6843 4326 6855 4378
rect 6855 4326 6869 4378
rect 6893 4326 6907 4378
rect 6907 4326 6919 4378
rect 6919 4326 6949 4378
rect 6973 4326 6983 4378
rect 6983 4326 7029 4378
rect 6733 4324 6789 4326
rect 6813 4324 6869 4326
rect 6893 4324 6949 4326
rect 6973 4324 7029 4326
rect 6733 3290 6789 3292
rect 6813 3290 6869 3292
rect 6893 3290 6949 3292
rect 6973 3290 7029 3292
rect 6733 3238 6779 3290
rect 6779 3238 6789 3290
rect 6813 3238 6843 3290
rect 6843 3238 6855 3290
rect 6855 3238 6869 3290
rect 6893 3238 6907 3290
rect 6907 3238 6919 3290
rect 6919 3238 6949 3290
rect 6973 3238 6983 3290
rect 6983 3238 7029 3290
rect 6733 3236 6789 3238
rect 6813 3236 6869 3238
rect 6893 3236 6949 3238
rect 6973 3236 7029 3238
rect 8120 4922 8176 4924
rect 8200 4922 8256 4924
rect 8280 4922 8336 4924
rect 8360 4922 8416 4924
rect 8120 4870 8166 4922
rect 8166 4870 8176 4922
rect 8200 4870 8230 4922
rect 8230 4870 8242 4922
rect 8242 4870 8256 4922
rect 8280 4870 8294 4922
rect 8294 4870 8306 4922
rect 8306 4870 8336 4922
rect 8360 4870 8370 4922
rect 8370 4870 8416 4922
rect 8120 4868 8176 4870
rect 8200 4868 8256 4870
rect 8280 4868 8336 4870
rect 8360 4868 8416 4870
rect 8780 6554 8836 6556
rect 8860 6554 8916 6556
rect 8940 6554 8996 6556
rect 9020 6554 9076 6556
rect 8780 6502 8826 6554
rect 8826 6502 8836 6554
rect 8860 6502 8890 6554
rect 8890 6502 8902 6554
rect 8902 6502 8916 6554
rect 8940 6502 8954 6554
rect 8954 6502 8966 6554
rect 8966 6502 8996 6554
rect 9020 6502 9030 6554
rect 9030 6502 9076 6554
rect 8780 6500 8836 6502
rect 8860 6500 8916 6502
rect 8940 6500 8996 6502
rect 9020 6500 9076 6502
rect 8780 5466 8836 5468
rect 8860 5466 8916 5468
rect 8940 5466 8996 5468
rect 9020 5466 9076 5468
rect 8780 5414 8826 5466
rect 8826 5414 8836 5466
rect 8860 5414 8890 5466
rect 8890 5414 8902 5466
rect 8902 5414 8916 5466
rect 8940 5414 8954 5466
rect 8954 5414 8966 5466
rect 8966 5414 8996 5466
rect 9020 5414 9030 5466
rect 9030 5414 9076 5466
rect 8780 5412 8836 5414
rect 8860 5412 8916 5414
rect 8940 5412 8996 5414
rect 9020 5412 9076 5414
rect 8758 5228 8814 5264
rect 8758 5208 8760 5228
rect 8760 5208 8812 5228
rect 8812 5208 8814 5228
rect 8780 4378 8836 4380
rect 8860 4378 8916 4380
rect 8940 4378 8996 4380
rect 9020 4378 9076 4380
rect 8780 4326 8826 4378
rect 8826 4326 8836 4378
rect 8860 4326 8890 4378
rect 8890 4326 8902 4378
rect 8902 4326 8916 4378
rect 8940 4326 8954 4378
rect 8954 4326 8966 4378
rect 8966 4326 8996 4378
rect 9020 4326 9030 4378
rect 9030 4326 9076 4378
rect 8780 4324 8836 4326
rect 8860 4324 8916 4326
rect 8940 4324 8996 4326
rect 9020 4324 9076 4326
rect 8120 3834 8176 3836
rect 8200 3834 8256 3836
rect 8280 3834 8336 3836
rect 8360 3834 8416 3836
rect 8120 3782 8166 3834
rect 8166 3782 8176 3834
rect 8200 3782 8230 3834
rect 8230 3782 8242 3834
rect 8242 3782 8256 3834
rect 8280 3782 8294 3834
rect 8294 3782 8306 3834
rect 8306 3782 8336 3834
rect 8360 3782 8370 3834
rect 8370 3782 8416 3834
rect 8120 3780 8176 3782
rect 8200 3780 8256 3782
rect 8280 3780 8336 3782
rect 8360 3780 8416 3782
rect 8780 3290 8836 3292
rect 8860 3290 8916 3292
rect 8940 3290 8996 3292
rect 9020 3290 9076 3292
rect 8780 3238 8826 3290
rect 8826 3238 8836 3290
rect 8860 3238 8890 3290
rect 8890 3238 8902 3290
rect 8902 3238 8916 3290
rect 8940 3238 8954 3290
rect 8954 3238 8966 3290
rect 8966 3238 8996 3290
rect 9020 3238 9030 3290
rect 9030 3238 9076 3290
rect 8780 3236 8836 3238
rect 8860 3236 8916 3238
rect 8940 3236 8996 3238
rect 9020 3236 9076 3238
rect 8120 2746 8176 2748
rect 8200 2746 8256 2748
rect 8280 2746 8336 2748
rect 8360 2746 8416 2748
rect 8120 2694 8166 2746
rect 8166 2694 8176 2746
rect 8200 2694 8230 2746
rect 8230 2694 8242 2746
rect 8242 2694 8256 2746
rect 8280 2694 8294 2746
rect 8294 2694 8306 2746
rect 8306 2694 8336 2746
rect 8360 2694 8370 2746
rect 8370 2694 8416 2746
rect 8120 2692 8176 2694
rect 8200 2692 8256 2694
rect 8280 2692 8336 2694
rect 8360 2692 8416 2694
rect 2639 2202 2695 2204
rect 2719 2202 2775 2204
rect 2799 2202 2855 2204
rect 2879 2202 2935 2204
rect 2639 2150 2685 2202
rect 2685 2150 2695 2202
rect 2719 2150 2749 2202
rect 2749 2150 2761 2202
rect 2761 2150 2775 2202
rect 2799 2150 2813 2202
rect 2813 2150 2825 2202
rect 2825 2150 2855 2202
rect 2879 2150 2889 2202
rect 2889 2150 2935 2202
rect 2639 2148 2695 2150
rect 2719 2148 2775 2150
rect 2799 2148 2855 2150
rect 2879 2148 2935 2150
rect 4686 2202 4742 2204
rect 4766 2202 4822 2204
rect 4846 2202 4902 2204
rect 4926 2202 4982 2204
rect 4686 2150 4732 2202
rect 4732 2150 4742 2202
rect 4766 2150 4796 2202
rect 4796 2150 4808 2202
rect 4808 2150 4822 2202
rect 4846 2150 4860 2202
rect 4860 2150 4872 2202
rect 4872 2150 4902 2202
rect 4926 2150 4936 2202
rect 4936 2150 4982 2202
rect 4686 2148 4742 2150
rect 4766 2148 4822 2150
rect 4846 2148 4902 2150
rect 4926 2148 4982 2150
rect 6733 2202 6789 2204
rect 6813 2202 6869 2204
rect 6893 2202 6949 2204
rect 6973 2202 7029 2204
rect 6733 2150 6779 2202
rect 6779 2150 6789 2202
rect 6813 2150 6843 2202
rect 6843 2150 6855 2202
rect 6855 2150 6869 2202
rect 6893 2150 6907 2202
rect 6907 2150 6919 2202
rect 6919 2150 6949 2202
rect 6973 2150 6983 2202
rect 6983 2150 7029 2202
rect 6733 2148 6789 2150
rect 6813 2148 6869 2150
rect 6893 2148 6949 2150
rect 6973 2148 7029 2150
rect 8780 2202 8836 2204
rect 8860 2202 8916 2204
rect 8940 2202 8996 2204
rect 9020 2202 9076 2204
rect 8780 2150 8826 2202
rect 8826 2150 8836 2202
rect 8860 2150 8890 2202
rect 8890 2150 8902 2202
rect 8902 2150 8916 2202
rect 8940 2150 8954 2202
rect 8954 2150 8966 2202
rect 8966 2150 8996 2202
rect 9020 2150 9030 2202
rect 9030 2150 9076 2202
rect 8780 2148 8836 2150
rect 8860 2148 8916 2150
rect 8940 2148 8996 2150
rect 9020 2148 9076 2150
<< metal3 >>
rect 1969 10368 2285 10369
rect 1969 10304 1975 10368
rect 2039 10304 2055 10368
rect 2119 10304 2135 10368
rect 2199 10304 2215 10368
rect 2279 10304 2285 10368
rect 1969 10303 2285 10304
rect 4016 10368 4332 10369
rect 4016 10304 4022 10368
rect 4086 10304 4102 10368
rect 4166 10304 4182 10368
rect 4246 10304 4262 10368
rect 4326 10304 4332 10368
rect 4016 10303 4332 10304
rect 6063 10368 6379 10369
rect 6063 10304 6069 10368
rect 6133 10304 6149 10368
rect 6213 10304 6229 10368
rect 6293 10304 6309 10368
rect 6373 10304 6379 10368
rect 6063 10303 6379 10304
rect 8110 10368 8426 10369
rect 8110 10304 8116 10368
rect 8180 10304 8196 10368
rect 8260 10304 8276 10368
rect 8340 10304 8356 10368
rect 8420 10304 8426 10368
rect 8110 10303 8426 10304
rect 2629 9824 2945 9825
rect 2629 9760 2635 9824
rect 2699 9760 2715 9824
rect 2779 9760 2795 9824
rect 2859 9760 2875 9824
rect 2939 9760 2945 9824
rect 2629 9759 2945 9760
rect 4676 9824 4992 9825
rect 4676 9760 4682 9824
rect 4746 9760 4762 9824
rect 4826 9760 4842 9824
rect 4906 9760 4922 9824
rect 4986 9760 4992 9824
rect 4676 9759 4992 9760
rect 6723 9824 7039 9825
rect 6723 9760 6729 9824
rect 6793 9760 6809 9824
rect 6873 9760 6889 9824
rect 6953 9760 6969 9824
rect 7033 9760 7039 9824
rect 6723 9759 7039 9760
rect 8770 9824 9086 9825
rect 8770 9760 8776 9824
rect 8840 9760 8856 9824
rect 8920 9760 8936 9824
rect 9000 9760 9016 9824
rect 9080 9760 9086 9824
rect 8770 9759 9086 9760
rect 0 9618 800 9648
rect 4429 9618 4495 9621
rect 0 9616 4495 9618
rect 0 9560 4434 9616
rect 4490 9560 4495 9616
rect 0 9558 4495 9560
rect 0 9528 800 9558
rect 4429 9555 4495 9558
rect 1969 9280 2285 9281
rect 1969 9216 1975 9280
rect 2039 9216 2055 9280
rect 2119 9216 2135 9280
rect 2199 9216 2215 9280
rect 2279 9216 2285 9280
rect 1969 9215 2285 9216
rect 4016 9280 4332 9281
rect 4016 9216 4022 9280
rect 4086 9216 4102 9280
rect 4166 9216 4182 9280
rect 4246 9216 4262 9280
rect 4326 9216 4332 9280
rect 4016 9215 4332 9216
rect 6063 9280 6379 9281
rect 6063 9216 6069 9280
rect 6133 9216 6149 9280
rect 6213 9216 6229 9280
rect 6293 9216 6309 9280
rect 6373 9216 6379 9280
rect 6063 9215 6379 9216
rect 8110 9280 8426 9281
rect 8110 9216 8116 9280
rect 8180 9216 8196 9280
rect 8260 9216 8276 9280
rect 8340 9216 8356 9280
rect 8420 9216 8426 9280
rect 8110 9215 8426 9216
rect 1577 8938 1643 8941
rect 3969 8938 4035 8941
rect 1577 8936 4035 8938
rect 1577 8880 1582 8936
rect 1638 8880 3974 8936
rect 4030 8880 4035 8936
rect 1577 8878 4035 8880
rect 1577 8875 1643 8878
rect 3969 8875 4035 8878
rect 6177 8938 6243 8941
rect 7557 8938 7623 8941
rect 6177 8936 7623 8938
rect 6177 8880 6182 8936
rect 6238 8880 7562 8936
rect 7618 8880 7623 8936
rect 6177 8878 7623 8880
rect 6177 8875 6243 8878
rect 7557 8875 7623 8878
rect 2629 8736 2945 8737
rect 2629 8672 2635 8736
rect 2699 8672 2715 8736
rect 2779 8672 2795 8736
rect 2859 8672 2875 8736
rect 2939 8672 2945 8736
rect 2629 8671 2945 8672
rect 4676 8736 4992 8737
rect 4676 8672 4682 8736
rect 4746 8672 4762 8736
rect 4826 8672 4842 8736
rect 4906 8672 4922 8736
rect 4986 8672 4992 8736
rect 4676 8671 4992 8672
rect 6723 8736 7039 8737
rect 6723 8672 6729 8736
rect 6793 8672 6809 8736
rect 6873 8672 6889 8736
rect 6953 8672 6969 8736
rect 7033 8672 7039 8736
rect 6723 8671 7039 8672
rect 8770 8736 9086 8737
rect 8770 8672 8776 8736
rect 8840 8672 8856 8736
rect 8920 8672 8936 8736
rect 9000 8672 9016 8736
rect 9080 8672 9086 8736
rect 8770 8671 9086 8672
rect 1853 8394 1919 8397
rect 3601 8394 3667 8397
rect 1853 8392 3667 8394
rect 1853 8336 1858 8392
rect 1914 8336 3606 8392
rect 3662 8336 3667 8392
rect 1853 8334 3667 8336
rect 1853 8331 1919 8334
rect 3601 8331 3667 8334
rect 1969 8192 2285 8193
rect 1969 8128 1975 8192
rect 2039 8128 2055 8192
rect 2119 8128 2135 8192
rect 2199 8128 2215 8192
rect 2279 8128 2285 8192
rect 1969 8127 2285 8128
rect 4016 8192 4332 8193
rect 4016 8128 4022 8192
rect 4086 8128 4102 8192
rect 4166 8128 4182 8192
rect 4246 8128 4262 8192
rect 4326 8128 4332 8192
rect 4016 8127 4332 8128
rect 6063 8192 6379 8193
rect 6063 8128 6069 8192
rect 6133 8128 6149 8192
rect 6213 8128 6229 8192
rect 6293 8128 6309 8192
rect 6373 8128 6379 8192
rect 6063 8127 6379 8128
rect 8110 8192 8426 8193
rect 8110 8128 8116 8192
rect 8180 8128 8196 8192
rect 8260 8128 8276 8192
rect 8340 8128 8356 8192
rect 8420 8128 8426 8192
rect 8110 8127 8426 8128
rect 2957 7986 3023 7989
rect 3325 7986 3391 7989
rect 2957 7984 3391 7986
rect 2957 7928 2962 7984
rect 3018 7928 3330 7984
rect 3386 7928 3391 7984
rect 2957 7926 3391 7928
rect 2957 7923 3023 7926
rect 3325 7923 3391 7926
rect 2313 7850 2379 7853
rect 3601 7850 3667 7853
rect 2313 7848 3667 7850
rect 2313 7792 2318 7848
rect 2374 7792 3606 7848
rect 3662 7792 3667 7848
rect 2313 7790 3667 7792
rect 2313 7787 2379 7790
rect 3601 7787 3667 7790
rect 2629 7648 2945 7649
rect 2629 7584 2635 7648
rect 2699 7584 2715 7648
rect 2779 7584 2795 7648
rect 2859 7584 2875 7648
rect 2939 7584 2945 7648
rect 2629 7583 2945 7584
rect 4676 7648 4992 7649
rect 4676 7584 4682 7648
rect 4746 7584 4762 7648
rect 4826 7584 4842 7648
rect 4906 7584 4922 7648
rect 4986 7584 4992 7648
rect 4676 7583 4992 7584
rect 6723 7648 7039 7649
rect 6723 7584 6729 7648
rect 6793 7584 6809 7648
rect 6873 7584 6889 7648
rect 6953 7584 6969 7648
rect 7033 7584 7039 7648
rect 6723 7583 7039 7584
rect 8770 7648 9086 7649
rect 8770 7584 8776 7648
rect 8840 7584 8856 7648
rect 8920 7584 8936 7648
rect 9000 7584 9016 7648
rect 9080 7584 9086 7648
rect 8770 7583 9086 7584
rect 5349 7578 5415 7581
rect 5349 7576 6562 7578
rect 5349 7520 5354 7576
rect 5410 7520 6562 7576
rect 5349 7518 6562 7520
rect 5349 7515 5415 7518
rect 4981 7442 5047 7445
rect 5758 7442 5764 7444
rect 4981 7440 5764 7442
rect 4981 7384 4986 7440
rect 5042 7384 5764 7440
rect 4981 7382 5764 7384
rect 4981 7379 5047 7382
rect 5758 7380 5764 7382
rect 5828 7442 5834 7444
rect 5993 7442 6059 7445
rect 5828 7440 6059 7442
rect 5828 7384 5998 7440
rect 6054 7384 6059 7440
rect 5828 7382 6059 7384
rect 6502 7442 6562 7518
rect 7281 7442 7347 7445
rect 6502 7440 7347 7442
rect 6502 7384 7286 7440
rect 7342 7384 7347 7440
rect 6502 7382 7347 7384
rect 5828 7380 5834 7382
rect 5993 7379 6059 7382
rect 7281 7379 7347 7382
rect 1969 7104 2285 7105
rect 1969 7040 1975 7104
rect 2039 7040 2055 7104
rect 2119 7040 2135 7104
rect 2199 7040 2215 7104
rect 2279 7040 2285 7104
rect 1969 7039 2285 7040
rect 4016 7104 4332 7105
rect 4016 7040 4022 7104
rect 4086 7040 4102 7104
rect 4166 7040 4182 7104
rect 4246 7040 4262 7104
rect 4326 7040 4332 7104
rect 4016 7039 4332 7040
rect 6063 7104 6379 7105
rect 6063 7040 6069 7104
rect 6133 7040 6149 7104
rect 6213 7040 6229 7104
rect 6293 7040 6309 7104
rect 6373 7040 6379 7104
rect 6063 7039 6379 7040
rect 8110 7104 8426 7105
rect 8110 7040 8116 7104
rect 8180 7040 8196 7104
rect 8260 7040 8276 7104
rect 8340 7040 8356 7104
rect 8420 7040 8426 7104
rect 8110 7039 8426 7040
rect 4981 7034 5047 7037
rect 4981 7032 5826 7034
rect 4981 6976 4986 7032
rect 5042 6976 5826 7032
rect 4981 6974 5826 6976
rect 4981 6971 5047 6974
rect 1945 6898 2011 6901
rect 4889 6898 4955 6901
rect 1945 6896 4955 6898
rect 1945 6840 1950 6896
rect 2006 6840 4894 6896
rect 4950 6840 4955 6896
rect 1945 6838 4955 6840
rect 5766 6898 5826 6974
rect 6177 6898 6243 6901
rect 5766 6896 6243 6898
rect 5766 6840 6182 6896
rect 6238 6840 6243 6896
rect 5766 6838 6243 6840
rect 1945 6835 2011 6838
rect 4889 6835 4955 6838
rect 6177 6835 6243 6838
rect 3509 6762 3575 6765
rect 3785 6762 3851 6765
rect 3509 6760 3851 6762
rect 3509 6704 3514 6760
rect 3570 6704 3790 6760
rect 3846 6704 3851 6760
rect 3509 6702 3851 6704
rect 3509 6699 3575 6702
rect 3785 6699 3851 6702
rect 4061 6762 4127 6765
rect 6821 6762 6887 6765
rect 4061 6760 6887 6762
rect 4061 6704 4066 6760
rect 4122 6704 6826 6760
rect 6882 6704 6887 6760
rect 4061 6702 6887 6704
rect 4061 6699 4127 6702
rect 6821 6699 6887 6702
rect 3233 6626 3299 6629
rect 3693 6626 3759 6629
rect 3233 6624 3759 6626
rect 3233 6568 3238 6624
rect 3294 6568 3698 6624
rect 3754 6568 3759 6624
rect 3233 6566 3759 6568
rect 3233 6563 3299 6566
rect 3693 6563 3759 6566
rect 2629 6560 2945 6561
rect 2629 6496 2635 6560
rect 2699 6496 2715 6560
rect 2779 6496 2795 6560
rect 2859 6496 2875 6560
rect 2939 6496 2945 6560
rect 2629 6495 2945 6496
rect 4676 6560 4992 6561
rect 4676 6496 4682 6560
rect 4746 6496 4762 6560
rect 4826 6496 4842 6560
rect 4906 6496 4922 6560
rect 4986 6496 4992 6560
rect 4676 6495 4992 6496
rect 6723 6560 7039 6561
rect 6723 6496 6729 6560
rect 6793 6496 6809 6560
rect 6873 6496 6889 6560
rect 6953 6496 6969 6560
rect 7033 6496 7039 6560
rect 6723 6495 7039 6496
rect 8770 6560 9086 6561
rect 8770 6496 8776 6560
rect 8840 6496 8856 6560
rect 8920 6496 8936 6560
rect 9000 6496 9016 6560
rect 9080 6496 9086 6560
rect 8770 6495 9086 6496
rect 3233 6490 3299 6493
rect 3969 6490 4035 6493
rect 3233 6488 4035 6490
rect 3233 6432 3238 6488
rect 3294 6432 3974 6488
rect 4030 6432 4035 6488
rect 3233 6430 4035 6432
rect 3233 6427 3299 6430
rect 3969 6427 4035 6430
rect 0 6218 800 6248
rect 1301 6218 1367 6221
rect 0 6216 1367 6218
rect 0 6160 1306 6216
rect 1362 6160 1367 6216
rect 0 6158 1367 6160
rect 0 6128 800 6158
rect 1301 6155 1367 6158
rect 1577 6218 1643 6221
rect 3969 6218 4035 6221
rect 1577 6216 4035 6218
rect 1577 6160 1582 6216
rect 1638 6160 3974 6216
rect 4030 6160 4035 6216
rect 1577 6158 4035 6160
rect 1577 6155 1643 6158
rect 3969 6155 4035 6158
rect 6361 6218 6427 6221
rect 6729 6218 6795 6221
rect 6361 6216 6795 6218
rect 6361 6160 6366 6216
rect 6422 6160 6734 6216
rect 6790 6160 6795 6216
rect 6361 6158 6795 6160
rect 6361 6155 6427 6158
rect 6729 6155 6795 6158
rect 1969 6016 2285 6017
rect 1969 5952 1975 6016
rect 2039 5952 2055 6016
rect 2119 5952 2135 6016
rect 2199 5952 2215 6016
rect 2279 5952 2285 6016
rect 1969 5951 2285 5952
rect 4016 6016 4332 6017
rect 4016 5952 4022 6016
rect 4086 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4332 6016
rect 4016 5951 4332 5952
rect 6063 6016 6379 6017
rect 6063 5952 6069 6016
rect 6133 5952 6149 6016
rect 6213 5952 6229 6016
rect 6293 5952 6309 6016
rect 6373 5952 6379 6016
rect 6063 5951 6379 5952
rect 8110 6016 8426 6017
rect 8110 5952 8116 6016
rect 8180 5952 8196 6016
rect 8260 5952 8276 6016
rect 8340 5952 8356 6016
rect 8420 5952 8426 6016
rect 8110 5951 8426 5952
rect 2865 5674 2931 5677
rect 3325 5674 3391 5677
rect 2865 5672 3391 5674
rect 2865 5616 2870 5672
rect 2926 5616 3330 5672
rect 3386 5616 3391 5672
rect 2865 5614 3391 5616
rect 2865 5611 2931 5614
rect 3325 5611 3391 5614
rect 5349 5674 5415 5677
rect 7465 5674 7531 5677
rect 5349 5672 7531 5674
rect 5349 5616 5354 5672
rect 5410 5616 7470 5672
rect 7526 5616 7531 5672
rect 5349 5614 7531 5616
rect 5349 5611 5415 5614
rect 7465 5611 7531 5614
rect 0 5538 800 5568
rect 0 5478 1042 5538
rect 0 5448 800 5478
rect 982 5266 1042 5478
rect 2629 5472 2945 5473
rect 2629 5408 2635 5472
rect 2699 5408 2715 5472
rect 2779 5408 2795 5472
rect 2859 5408 2875 5472
rect 2939 5408 2945 5472
rect 2629 5407 2945 5408
rect 4676 5472 4992 5473
rect 4676 5408 4682 5472
rect 4746 5408 4762 5472
rect 4826 5408 4842 5472
rect 4906 5408 4922 5472
rect 4986 5408 4992 5472
rect 4676 5407 4992 5408
rect 6723 5472 7039 5473
rect 6723 5408 6729 5472
rect 6793 5408 6809 5472
rect 6873 5408 6889 5472
rect 6953 5408 6969 5472
rect 7033 5408 7039 5472
rect 6723 5407 7039 5408
rect 8770 5472 9086 5473
rect 8770 5408 8776 5472
rect 8840 5408 8856 5472
rect 8920 5408 8936 5472
rect 9000 5408 9016 5472
rect 9080 5408 9086 5472
rect 8770 5407 9086 5408
rect 1761 5266 1827 5269
rect 982 5264 1827 5266
rect 982 5208 1766 5264
rect 1822 5208 1827 5264
rect 982 5206 1827 5208
rect 1761 5203 1827 5206
rect 6269 5266 6335 5269
rect 8753 5266 8819 5269
rect 6269 5264 8819 5266
rect 6269 5208 6274 5264
rect 6330 5208 8758 5264
rect 8814 5208 8819 5264
rect 6269 5206 8819 5208
rect 6269 5203 6335 5206
rect 8753 5203 8819 5206
rect 1969 4928 2285 4929
rect 1969 4864 1975 4928
rect 2039 4864 2055 4928
rect 2119 4864 2135 4928
rect 2199 4864 2215 4928
rect 2279 4864 2285 4928
rect 1969 4863 2285 4864
rect 4016 4928 4332 4929
rect 4016 4864 4022 4928
rect 4086 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4332 4928
rect 4016 4863 4332 4864
rect 6063 4928 6379 4929
rect 6063 4864 6069 4928
rect 6133 4864 6149 4928
rect 6213 4864 6229 4928
rect 6293 4864 6309 4928
rect 6373 4864 6379 4928
rect 6063 4863 6379 4864
rect 8110 4928 8426 4929
rect 8110 4864 8116 4928
rect 8180 4864 8196 4928
rect 8260 4864 8276 4928
rect 8340 4864 8356 4928
rect 8420 4864 8426 4928
rect 8110 4863 8426 4864
rect 5758 4660 5764 4724
rect 5828 4722 5834 4724
rect 6269 4722 6335 4725
rect 5828 4720 6335 4722
rect 5828 4664 6274 4720
rect 6330 4664 6335 4720
rect 5828 4662 6335 4664
rect 5828 4660 5834 4662
rect 6269 4659 6335 4662
rect 4429 4586 4495 4589
rect 5717 4586 5783 4589
rect 4429 4584 5783 4586
rect 4429 4528 4434 4584
rect 4490 4528 5722 4584
rect 5778 4528 5783 4584
rect 4429 4526 5783 4528
rect 4429 4523 4495 4526
rect 5717 4523 5783 4526
rect 2629 4384 2945 4385
rect 2629 4320 2635 4384
rect 2699 4320 2715 4384
rect 2779 4320 2795 4384
rect 2859 4320 2875 4384
rect 2939 4320 2945 4384
rect 2629 4319 2945 4320
rect 4676 4384 4992 4385
rect 4676 4320 4682 4384
rect 4746 4320 4762 4384
rect 4826 4320 4842 4384
rect 4906 4320 4922 4384
rect 4986 4320 4992 4384
rect 4676 4319 4992 4320
rect 6723 4384 7039 4385
rect 6723 4320 6729 4384
rect 6793 4320 6809 4384
rect 6873 4320 6889 4384
rect 6953 4320 6969 4384
rect 7033 4320 7039 4384
rect 6723 4319 7039 4320
rect 8770 4384 9086 4385
rect 8770 4320 8776 4384
rect 8840 4320 8856 4384
rect 8920 4320 8936 4384
rect 9000 4320 9016 4384
rect 9080 4320 9086 4384
rect 8770 4319 9086 4320
rect 2405 4042 2471 4045
rect 5625 4042 5691 4045
rect 2405 4040 5691 4042
rect 2405 3984 2410 4040
rect 2466 3984 5630 4040
rect 5686 3984 5691 4040
rect 2405 3982 5691 3984
rect 2405 3979 2471 3982
rect 5625 3979 5691 3982
rect 1969 3840 2285 3841
rect 1969 3776 1975 3840
rect 2039 3776 2055 3840
rect 2119 3776 2135 3840
rect 2199 3776 2215 3840
rect 2279 3776 2285 3840
rect 1969 3775 2285 3776
rect 4016 3840 4332 3841
rect 4016 3776 4022 3840
rect 4086 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4332 3840
rect 4016 3775 4332 3776
rect 6063 3840 6379 3841
rect 6063 3776 6069 3840
rect 6133 3776 6149 3840
rect 6213 3776 6229 3840
rect 6293 3776 6309 3840
rect 6373 3776 6379 3840
rect 6063 3775 6379 3776
rect 8110 3840 8426 3841
rect 8110 3776 8116 3840
rect 8180 3776 8196 3840
rect 8260 3776 8276 3840
rect 8340 3776 8356 3840
rect 8420 3776 8426 3840
rect 8110 3775 8426 3776
rect 4705 3498 4771 3501
rect 5533 3498 5599 3501
rect 4705 3496 5599 3498
rect 4705 3440 4710 3496
rect 4766 3440 5538 3496
rect 5594 3440 5599 3496
rect 4705 3438 5599 3440
rect 4705 3435 4771 3438
rect 5533 3435 5599 3438
rect 2629 3296 2945 3297
rect 2629 3232 2635 3296
rect 2699 3232 2715 3296
rect 2779 3232 2795 3296
rect 2859 3232 2875 3296
rect 2939 3232 2945 3296
rect 2629 3231 2945 3232
rect 4676 3296 4992 3297
rect 4676 3232 4682 3296
rect 4746 3232 4762 3296
rect 4826 3232 4842 3296
rect 4906 3232 4922 3296
rect 4986 3232 4992 3296
rect 4676 3231 4992 3232
rect 6723 3296 7039 3297
rect 6723 3232 6729 3296
rect 6793 3232 6809 3296
rect 6873 3232 6889 3296
rect 6953 3232 6969 3296
rect 7033 3232 7039 3296
rect 6723 3231 7039 3232
rect 8770 3296 9086 3297
rect 8770 3232 8776 3296
rect 8840 3232 8856 3296
rect 8920 3232 8936 3296
rect 9000 3232 9016 3296
rect 9080 3232 9086 3296
rect 8770 3231 9086 3232
rect 1969 2752 2285 2753
rect 1969 2688 1975 2752
rect 2039 2688 2055 2752
rect 2119 2688 2135 2752
rect 2199 2688 2215 2752
rect 2279 2688 2285 2752
rect 1969 2687 2285 2688
rect 4016 2752 4332 2753
rect 4016 2688 4022 2752
rect 4086 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4332 2752
rect 4016 2687 4332 2688
rect 6063 2752 6379 2753
rect 6063 2688 6069 2752
rect 6133 2688 6149 2752
rect 6213 2688 6229 2752
rect 6293 2688 6309 2752
rect 6373 2688 6379 2752
rect 6063 2687 6379 2688
rect 8110 2752 8426 2753
rect 8110 2688 8116 2752
rect 8180 2688 8196 2752
rect 8260 2688 8276 2752
rect 8340 2688 8356 2752
rect 8420 2688 8426 2752
rect 8110 2687 8426 2688
rect 2629 2208 2945 2209
rect 2629 2144 2635 2208
rect 2699 2144 2715 2208
rect 2779 2144 2795 2208
rect 2859 2144 2875 2208
rect 2939 2144 2945 2208
rect 2629 2143 2945 2144
rect 4676 2208 4992 2209
rect 4676 2144 4682 2208
rect 4746 2144 4762 2208
rect 4826 2144 4842 2208
rect 4906 2144 4922 2208
rect 4986 2144 4992 2208
rect 4676 2143 4992 2144
rect 6723 2208 7039 2209
rect 6723 2144 6729 2208
rect 6793 2144 6809 2208
rect 6873 2144 6889 2208
rect 6953 2144 6969 2208
rect 7033 2144 7039 2208
rect 6723 2143 7039 2144
rect 8770 2208 9086 2209
rect 8770 2144 8776 2208
rect 8840 2144 8856 2208
rect 8920 2144 8936 2208
rect 9000 2144 9016 2208
rect 9080 2144 9086 2208
rect 8770 2143 9086 2144
<< via3 >>
rect 1975 10364 2039 10368
rect 1975 10308 1979 10364
rect 1979 10308 2035 10364
rect 2035 10308 2039 10364
rect 1975 10304 2039 10308
rect 2055 10364 2119 10368
rect 2055 10308 2059 10364
rect 2059 10308 2115 10364
rect 2115 10308 2119 10364
rect 2055 10304 2119 10308
rect 2135 10364 2199 10368
rect 2135 10308 2139 10364
rect 2139 10308 2195 10364
rect 2195 10308 2199 10364
rect 2135 10304 2199 10308
rect 2215 10364 2279 10368
rect 2215 10308 2219 10364
rect 2219 10308 2275 10364
rect 2275 10308 2279 10364
rect 2215 10304 2279 10308
rect 4022 10364 4086 10368
rect 4022 10308 4026 10364
rect 4026 10308 4082 10364
rect 4082 10308 4086 10364
rect 4022 10304 4086 10308
rect 4102 10364 4166 10368
rect 4102 10308 4106 10364
rect 4106 10308 4162 10364
rect 4162 10308 4166 10364
rect 4102 10304 4166 10308
rect 4182 10364 4246 10368
rect 4182 10308 4186 10364
rect 4186 10308 4242 10364
rect 4242 10308 4246 10364
rect 4182 10304 4246 10308
rect 4262 10364 4326 10368
rect 4262 10308 4266 10364
rect 4266 10308 4322 10364
rect 4322 10308 4326 10364
rect 4262 10304 4326 10308
rect 6069 10364 6133 10368
rect 6069 10308 6073 10364
rect 6073 10308 6129 10364
rect 6129 10308 6133 10364
rect 6069 10304 6133 10308
rect 6149 10364 6213 10368
rect 6149 10308 6153 10364
rect 6153 10308 6209 10364
rect 6209 10308 6213 10364
rect 6149 10304 6213 10308
rect 6229 10364 6293 10368
rect 6229 10308 6233 10364
rect 6233 10308 6289 10364
rect 6289 10308 6293 10364
rect 6229 10304 6293 10308
rect 6309 10364 6373 10368
rect 6309 10308 6313 10364
rect 6313 10308 6369 10364
rect 6369 10308 6373 10364
rect 6309 10304 6373 10308
rect 8116 10364 8180 10368
rect 8116 10308 8120 10364
rect 8120 10308 8176 10364
rect 8176 10308 8180 10364
rect 8116 10304 8180 10308
rect 8196 10364 8260 10368
rect 8196 10308 8200 10364
rect 8200 10308 8256 10364
rect 8256 10308 8260 10364
rect 8196 10304 8260 10308
rect 8276 10364 8340 10368
rect 8276 10308 8280 10364
rect 8280 10308 8336 10364
rect 8336 10308 8340 10364
rect 8276 10304 8340 10308
rect 8356 10364 8420 10368
rect 8356 10308 8360 10364
rect 8360 10308 8416 10364
rect 8416 10308 8420 10364
rect 8356 10304 8420 10308
rect 2635 9820 2699 9824
rect 2635 9764 2639 9820
rect 2639 9764 2695 9820
rect 2695 9764 2699 9820
rect 2635 9760 2699 9764
rect 2715 9820 2779 9824
rect 2715 9764 2719 9820
rect 2719 9764 2775 9820
rect 2775 9764 2779 9820
rect 2715 9760 2779 9764
rect 2795 9820 2859 9824
rect 2795 9764 2799 9820
rect 2799 9764 2855 9820
rect 2855 9764 2859 9820
rect 2795 9760 2859 9764
rect 2875 9820 2939 9824
rect 2875 9764 2879 9820
rect 2879 9764 2935 9820
rect 2935 9764 2939 9820
rect 2875 9760 2939 9764
rect 4682 9820 4746 9824
rect 4682 9764 4686 9820
rect 4686 9764 4742 9820
rect 4742 9764 4746 9820
rect 4682 9760 4746 9764
rect 4762 9820 4826 9824
rect 4762 9764 4766 9820
rect 4766 9764 4822 9820
rect 4822 9764 4826 9820
rect 4762 9760 4826 9764
rect 4842 9820 4906 9824
rect 4842 9764 4846 9820
rect 4846 9764 4902 9820
rect 4902 9764 4906 9820
rect 4842 9760 4906 9764
rect 4922 9820 4986 9824
rect 4922 9764 4926 9820
rect 4926 9764 4982 9820
rect 4982 9764 4986 9820
rect 4922 9760 4986 9764
rect 6729 9820 6793 9824
rect 6729 9764 6733 9820
rect 6733 9764 6789 9820
rect 6789 9764 6793 9820
rect 6729 9760 6793 9764
rect 6809 9820 6873 9824
rect 6809 9764 6813 9820
rect 6813 9764 6869 9820
rect 6869 9764 6873 9820
rect 6809 9760 6873 9764
rect 6889 9820 6953 9824
rect 6889 9764 6893 9820
rect 6893 9764 6949 9820
rect 6949 9764 6953 9820
rect 6889 9760 6953 9764
rect 6969 9820 7033 9824
rect 6969 9764 6973 9820
rect 6973 9764 7029 9820
rect 7029 9764 7033 9820
rect 6969 9760 7033 9764
rect 8776 9820 8840 9824
rect 8776 9764 8780 9820
rect 8780 9764 8836 9820
rect 8836 9764 8840 9820
rect 8776 9760 8840 9764
rect 8856 9820 8920 9824
rect 8856 9764 8860 9820
rect 8860 9764 8916 9820
rect 8916 9764 8920 9820
rect 8856 9760 8920 9764
rect 8936 9820 9000 9824
rect 8936 9764 8940 9820
rect 8940 9764 8996 9820
rect 8996 9764 9000 9820
rect 8936 9760 9000 9764
rect 9016 9820 9080 9824
rect 9016 9764 9020 9820
rect 9020 9764 9076 9820
rect 9076 9764 9080 9820
rect 9016 9760 9080 9764
rect 1975 9276 2039 9280
rect 1975 9220 1979 9276
rect 1979 9220 2035 9276
rect 2035 9220 2039 9276
rect 1975 9216 2039 9220
rect 2055 9276 2119 9280
rect 2055 9220 2059 9276
rect 2059 9220 2115 9276
rect 2115 9220 2119 9276
rect 2055 9216 2119 9220
rect 2135 9276 2199 9280
rect 2135 9220 2139 9276
rect 2139 9220 2195 9276
rect 2195 9220 2199 9276
rect 2135 9216 2199 9220
rect 2215 9276 2279 9280
rect 2215 9220 2219 9276
rect 2219 9220 2275 9276
rect 2275 9220 2279 9276
rect 2215 9216 2279 9220
rect 4022 9276 4086 9280
rect 4022 9220 4026 9276
rect 4026 9220 4082 9276
rect 4082 9220 4086 9276
rect 4022 9216 4086 9220
rect 4102 9276 4166 9280
rect 4102 9220 4106 9276
rect 4106 9220 4162 9276
rect 4162 9220 4166 9276
rect 4102 9216 4166 9220
rect 4182 9276 4246 9280
rect 4182 9220 4186 9276
rect 4186 9220 4242 9276
rect 4242 9220 4246 9276
rect 4182 9216 4246 9220
rect 4262 9276 4326 9280
rect 4262 9220 4266 9276
rect 4266 9220 4322 9276
rect 4322 9220 4326 9276
rect 4262 9216 4326 9220
rect 6069 9276 6133 9280
rect 6069 9220 6073 9276
rect 6073 9220 6129 9276
rect 6129 9220 6133 9276
rect 6069 9216 6133 9220
rect 6149 9276 6213 9280
rect 6149 9220 6153 9276
rect 6153 9220 6209 9276
rect 6209 9220 6213 9276
rect 6149 9216 6213 9220
rect 6229 9276 6293 9280
rect 6229 9220 6233 9276
rect 6233 9220 6289 9276
rect 6289 9220 6293 9276
rect 6229 9216 6293 9220
rect 6309 9276 6373 9280
rect 6309 9220 6313 9276
rect 6313 9220 6369 9276
rect 6369 9220 6373 9276
rect 6309 9216 6373 9220
rect 8116 9276 8180 9280
rect 8116 9220 8120 9276
rect 8120 9220 8176 9276
rect 8176 9220 8180 9276
rect 8116 9216 8180 9220
rect 8196 9276 8260 9280
rect 8196 9220 8200 9276
rect 8200 9220 8256 9276
rect 8256 9220 8260 9276
rect 8196 9216 8260 9220
rect 8276 9276 8340 9280
rect 8276 9220 8280 9276
rect 8280 9220 8336 9276
rect 8336 9220 8340 9276
rect 8276 9216 8340 9220
rect 8356 9276 8420 9280
rect 8356 9220 8360 9276
rect 8360 9220 8416 9276
rect 8416 9220 8420 9276
rect 8356 9216 8420 9220
rect 2635 8732 2699 8736
rect 2635 8676 2639 8732
rect 2639 8676 2695 8732
rect 2695 8676 2699 8732
rect 2635 8672 2699 8676
rect 2715 8732 2779 8736
rect 2715 8676 2719 8732
rect 2719 8676 2775 8732
rect 2775 8676 2779 8732
rect 2715 8672 2779 8676
rect 2795 8732 2859 8736
rect 2795 8676 2799 8732
rect 2799 8676 2855 8732
rect 2855 8676 2859 8732
rect 2795 8672 2859 8676
rect 2875 8732 2939 8736
rect 2875 8676 2879 8732
rect 2879 8676 2935 8732
rect 2935 8676 2939 8732
rect 2875 8672 2939 8676
rect 4682 8732 4746 8736
rect 4682 8676 4686 8732
rect 4686 8676 4742 8732
rect 4742 8676 4746 8732
rect 4682 8672 4746 8676
rect 4762 8732 4826 8736
rect 4762 8676 4766 8732
rect 4766 8676 4822 8732
rect 4822 8676 4826 8732
rect 4762 8672 4826 8676
rect 4842 8732 4906 8736
rect 4842 8676 4846 8732
rect 4846 8676 4902 8732
rect 4902 8676 4906 8732
rect 4842 8672 4906 8676
rect 4922 8732 4986 8736
rect 4922 8676 4926 8732
rect 4926 8676 4982 8732
rect 4982 8676 4986 8732
rect 4922 8672 4986 8676
rect 6729 8732 6793 8736
rect 6729 8676 6733 8732
rect 6733 8676 6789 8732
rect 6789 8676 6793 8732
rect 6729 8672 6793 8676
rect 6809 8732 6873 8736
rect 6809 8676 6813 8732
rect 6813 8676 6869 8732
rect 6869 8676 6873 8732
rect 6809 8672 6873 8676
rect 6889 8732 6953 8736
rect 6889 8676 6893 8732
rect 6893 8676 6949 8732
rect 6949 8676 6953 8732
rect 6889 8672 6953 8676
rect 6969 8732 7033 8736
rect 6969 8676 6973 8732
rect 6973 8676 7029 8732
rect 7029 8676 7033 8732
rect 6969 8672 7033 8676
rect 8776 8732 8840 8736
rect 8776 8676 8780 8732
rect 8780 8676 8836 8732
rect 8836 8676 8840 8732
rect 8776 8672 8840 8676
rect 8856 8732 8920 8736
rect 8856 8676 8860 8732
rect 8860 8676 8916 8732
rect 8916 8676 8920 8732
rect 8856 8672 8920 8676
rect 8936 8732 9000 8736
rect 8936 8676 8940 8732
rect 8940 8676 8996 8732
rect 8996 8676 9000 8732
rect 8936 8672 9000 8676
rect 9016 8732 9080 8736
rect 9016 8676 9020 8732
rect 9020 8676 9076 8732
rect 9076 8676 9080 8732
rect 9016 8672 9080 8676
rect 1975 8188 2039 8192
rect 1975 8132 1979 8188
rect 1979 8132 2035 8188
rect 2035 8132 2039 8188
rect 1975 8128 2039 8132
rect 2055 8188 2119 8192
rect 2055 8132 2059 8188
rect 2059 8132 2115 8188
rect 2115 8132 2119 8188
rect 2055 8128 2119 8132
rect 2135 8188 2199 8192
rect 2135 8132 2139 8188
rect 2139 8132 2195 8188
rect 2195 8132 2199 8188
rect 2135 8128 2199 8132
rect 2215 8188 2279 8192
rect 2215 8132 2219 8188
rect 2219 8132 2275 8188
rect 2275 8132 2279 8188
rect 2215 8128 2279 8132
rect 4022 8188 4086 8192
rect 4022 8132 4026 8188
rect 4026 8132 4082 8188
rect 4082 8132 4086 8188
rect 4022 8128 4086 8132
rect 4102 8188 4166 8192
rect 4102 8132 4106 8188
rect 4106 8132 4162 8188
rect 4162 8132 4166 8188
rect 4102 8128 4166 8132
rect 4182 8188 4246 8192
rect 4182 8132 4186 8188
rect 4186 8132 4242 8188
rect 4242 8132 4246 8188
rect 4182 8128 4246 8132
rect 4262 8188 4326 8192
rect 4262 8132 4266 8188
rect 4266 8132 4322 8188
rect 4322 8132 4326 8188
rect 4262 8128 4326 8132
rect 6069 8188 6133 8192
rect 6069 8132 6073 8188
rect 6073 8132 6129 8188
rect 6129 8132 6133 8188
rect 6069 8128 6133 8132
rect 6149 8188 6213 8192
rect 6149 8132 6153 8188
rect 6153 8132 6209 8188
rect 6209 8132 6213 8188
rect 6149 8128 6213 8132
rect 6229 8188 6293 8192
rect 6229 8132 6233 8188
rect 6233 8132 6289 8188
rect 6289 8132 6293 8188
rect 6229 8128 6293 8132
rect 6309 8188 6373 8192
rect 6309 8132 6313 8188
rect 6313 8132 6369 8188
rect 6369 8132 6373 8188
rect 6309 8128 6373 8132
rect 8116 8188 8180 8192
rect 8116 8132 8120 8188
rect 8120 8132 8176 8188
rect 8176 8132 8180 8188
rect 8116 8128 8180 8132
rect 8196 8188 8260 8192
rect 8196 8132 8200 8188
rect 8200 8132 8256 8188
rect 8256 8132 8260 8188
rect 8196 8128 8260 8132
rect 8276 8188 8340 8192
rect 8276 8132 8280 8188
rect 8280 8132 8336 8188
rect 8336 8132 8340 8188
rect 8276 8128 8340 8132
rect 8356 8188 8420 8192
rect 8356 8132 8360 8188
rect 8360 8132 8416 8188
rect 8416 8132 8420 8188
rect 8356 8128 8420 8132
rect 2635 7644 2699 7648
rect 2635 7588 2639 7644
rect 2639 7588 2695 7644
rect 2695 7588 2699 7644
rect 2635 7584 2699 7588
rect 2715 7644 2779 7648
rect 2715 7588 2719 7644
rect 2719 7588 2775 7644
rect 2775 7588 2779 7644
rect 2715 7584 2779 7588
rect 2795 7644 2859 7648
rect 2795 7588 2799 7644
rect 2799 7588 2855 7644
rect 2855 7588 2859 7644
rect 2795 7584 2859 7588
rect 2875 7644 2939 7648
rect 2875 7588 2879 7644
rect 2879 7588 2935 7644
rect 2935 7588 2939 7644
rect 2875 7584 2939 7588
rect 4682 7644 4746 7648
rect 4682 7588 4686 7644
rect 4686 7588 4742 7644
rect 4742 7588 4746 7644
rect 4682 7584 4746 7588
rect 4762 7644 4826 7648
rect 4762 7588 4766 7644
rect 4766 7588 4822 7644
rect 4822 7588 4826 7644
rect 4762 7584 4826 7588
rect 4842 7644 4906 7648
rect 4842 7588 4846 7644
rect 4846 7588 4902 7644
rect 4902 7588 4906 7644
rect 4842 7584 4906 7588
rect 4922 7644 4986 7648
rect 4922 7588 4926 7644
rect 4926 7588 4982 7644
rect 4982 7588 4986 7644
rect 4922 7584 4986 7588
rect 6729 7644 6793 7648
rect 6729 7588 6733 7644
rect 6733 7588 6789 7644
rect 6789 7588 6793 7644
rect 6729 7584 6793 7588
rect 6809 7644 6873 7648
rect 6809 7588 6813 7644
rect 6813 7588 6869 7644
rect 6869 7588 6873 7644
rect 6809 7584 6873 7588
rect 6889 7644 6953 7648
rect 6889 7588 6893 7644
rect 6893 7588 6949 7644
rect 6949 7588 6953 7644
rect 6889 7584 6953 7588
rect 6969 7644 7033 7648
rect 6969 7588 6973 7644
rect 6973 7588 7029 7644
rect 7029 7588 7033 7644
rect 6969 7584 7033 7588
rect 8776 7644 8840 7648
rect 8776 7588 8780 7644
rect 8780 7588 8836 7644
rect 8836 7588 8840 7644
rect 8776 7584 8840 7588
rect 8856 7644 8920 7648
rect 8856 7588 8860 7644
rect 8860 7588 8916 7644
rect 8916 7588 8920 7644
rect 8856 7584 8920 7588
rect 8936 7644 9000 7648
rect 8936 7588 8940 7644
rect 8940 7588 8996 7644
rect 8996 7588 9000 7644
rect 8936 7584 9000 7588
rect 9016 7644 9080 7648
rect 9016 7588 9020 7644
rect 9020 7588 9076 7644
rect 9076 7588 9080 7644
rect 9016 7584 9080 7588
rect 5764 7380 5828 7444
rect 1975 7100 2039 7104
rect 1975 7044 1979 7100
rect 1979 7044 2035 7100
rect 2035 7044 2039 7100
rect 1975 7040 2039 7044
rect 2055 7100 2119 7104
rect 2055 7044 2059 7100
rect 2059 7044 2115 7100
rect 2115 7044 2119 7100
rect 2055 7040 2119 7044
rect 2135 7100 2199 7104
rect 2135 7044 2139 7100
rect 2139 7044 2195 7100
rect 2195 7044 2199 7100
rect 2135 7040 2199 7044
rect 2215 7100 2279 7104
rect 2215 7044 2219 7100
rect 2219 7044 2275 7100
rect 2275 7044 2279 7100
rect 2215 7040 2279 7044
rect 4022 7100 4086 7104
rect 4022 7044 4026 7100
rect 4026 7044 4082 7100
rect 4082 7044 4086 7100
rect 4022 7040 4086 7044
rect 4102 7100 4166 7104
rect 4102 7044 4106 7100
rect 4106 7044 4162 7100
rect 4162 7044 4166 7100
rect 4102 7040 4166 7044
rect 4182 7100 4246 7104
rect 4182 7044 4186 7100
rect 4186 7044 4242 7100
rect 4242 7044 4246 7100
rect 4182 7040 4246 7044
rect 4262 7100 4326 7104
rect 4262 7044 4266 7100
rect 4266 7044 4322 7100
rect 4322 7044 4326 7100
rect 4262 7040 4326 7044
rect 6069 7100 6133 7104
rect 6069 7044 6073 7100
rect 6073 7044 6129 7100
rect 6129 7044 6133 7100
rect 6069 7040 6133 7044
rect 6149 7100 6213 7104
rect 6149 7044 6153 7100
rect 6153 7044 6209 7100
rect 6209 7044 6213 7100
rect 6149 7040 6213 7044
rect 6229 7100 6293 7104
rect 6229 7044 6233 7100
rect 6233 7044 6289 7100
rect 6289 7044 6293 7100
rect 6229 7040 6293 7044
rect 6309 7100 6373 7104
rect 6309 7044 6313 7100
rect 6313 7044 6369 7100
rect 6369 7044 6373 7100
rect 6309 7040 6373 7044
rect 8116 7100 8180 7104
rect 8116 7044 8120 7100
rect 8120 7044 8176 7100
rect 8176 7044 8180 7100
rect 8116 7040 8180 7044
rect 8196 7100 8260 7104
rect 8196 7044 8200 7100
rect 8200 7044 8256 7100
rect 8256 7044 8260 7100
rect 8196 7040 8260 7044
rect 8276 7100 8340 7104
rect 8276 7044 8280 7100
rect 8280 7044 8336 7100
rect 8336 7044 8340 7100
rect 8276 7040 8340 7044
rect 8356 7100 8420 7104
rect 8356 7044 8360 7100
rect 8360 7044 8416 7100
rect 8416 7044 8420 7100
rect 8356 7040 8420 7044
rect 2635 6556 2699 6560
rect 2635 6500 2639 6556
rect 2639 6500 2695 6556
rect 2695 6500 2699 6556
rect 2635 6496 2699 6500
rect 2715 6556 2779 6560
rect 2715 6500 2719 6556
rect 2719 6500 2775 6556
rect 2775 6500 2779 6556
rect 2715 6496 2779 6500
rect 2795 6556 2859 6560
rect 2795 6500 2799 6556
rect 2799 6500 2855 6556
rect 2855 6500 2859 6556
rect 2795 6496 2859 6500
rect 2875 6556 2939 6560
rect 2875 6500 2879 6556
rect 2879 6500 2935 6556
rect 2935 6500 2939 6556
rect 2875 6496 2939 6500
rect 4682 6556 4746 6560
rect 4682 6500 4686 6556
rect 4686 6500 4742 6556
rect 4742 6500 4746 6556
rect 4682 6496 4746 6500
rect 4762 6556 4826 6560
rect 4762 6500 4766 6556
rect 4766 6500 4822 6556
rect 4822 6500 4826 6556
rect 4762 6496 4826 6500
rect 4842 6556 4906 6560
rect 4842 6500 4846 6556
rect 4846 6500 4902 6556
rect 4902 6500 4906 6556
rect 4842 6496 4906 6500
rect 4922 6556 4986 6560
rect 4922 6500 4926 6556
rect 4926 6500 4982 6556
rect 4982 6500 4986 6556
rect 4922 6496 4986 6500
rect 6729 6556 6793 6560
rect 6729 6500 6733 6556
rect 6733 6500 6789 6556
rect 6789 6500 6793 6556
rect 6729 6496 6793 6500
rect 6809 6556 6873 6560
rect 6809 6500 6813 6556
rect 6813 6500 6869 6556
rect 6869 6500 6873 6556
rect 6809 6496 6873 6500
rect 6889 6556 6953 6560
rect 6889 6500 6893 6556
rect 6893 6500 6949 6556
rect 6949 6500 6953 6556
rect 6889 6496 6953 6500
rect 6969 6556 7033 6560
rect 6969 6500 6973 6556
rect 6973 6500 7029 6556
rect 7029 6500 7033 6556
rect 6969 6496 7033 6500
rect 8776 6556 8840 6560
rect 8776 6500 8780 6556
rect 8780 6500 8836 6556
rect 8836 6500 8840 6556
rect 8776 6496 8840 6500
rect 8856 6556 8920 6560
rect 8856 6500 8860 6556
rect 8860 6500 8916 6556
rect 8916 6500 8920 6556
rect 8856 6496 8920 6500
rect 8936 6556 9000 6560
rect 8936 6500 8940 6556
rect 8940 6500 8996 6556
rect 8996 6500 9000 6556
rect 8936 6496 9000 6500
rect 9016 6556 9080 6560
rect 9016 6500 9020 6556
rect 9020 6500 9076 6556
rect 9076 6500 9080 6556
rect 9016 6496 9080 6500
rect 1975 6012 2039 6016
rect 1975 5956 1979 6012
rect 1979 5956 2035 6012
rect 2035 5956 2039 6012
rect 1975 5952 2039 5956
rect 2055 6012 2119 6016
rect 2055 5956 2059 6012
rect 2059 5956 2115 6012
rect 2115 5956 2119 6012
rect 2055 5952 2119 5956
rect 2135 6012 2199 6016
rect 2135 5956 2139 6012
rect 2139 5956 2195 6012
rect 2195 5956 2199 6012
rect 2135 5952 2199 5956
rect 2215 6012 2279 6016
rect 2215 5956 2219 6012
rect 2219 5956 2275 6012
rect 2275 5956 2279 6012
rect 2215 5952 2279 5956
rect 4022 6012 4086 6016
rect 4022 5956 4026 6012
rect 4026 5956 4082 6012
rect 4082 5956 4086 6012
rect 4022 5952 4086 5956
rect 4102 6012 4166 6016
rect 4102 5956 4106 6012
rect 4106 5956 4162 6012
rect 4162 5956 4166 6012
rect 4102 5952 4166 5956
rect 4182 6012 4246 6016
rect 4182 5956 4186 6012
rect 4186 5956 4242 6012
rect 4242 5956 4246 6012
rect 4182 5952 4246 5956
rect 4262 6012 4326 6016
rect 4262 5956 4266 6012
rect 4266 5956 4322 6012
rect 4322 5956 4326 6012
rect 4262 5952 4326 5956
rect 6069 6012 6133 6016
rect 6069 5956 6073 6012
rect 6073 5956 6129 6012
rect 6129 5956 6133 6012
rect 6069 5952 6133 5956
rect 6149 6012 6213 6016
rect 6149 5956 6153 6012
rect 6153 5956 6209 6012
rect 6209 5956 6213 6012
rect 6149 5952 6213 5956
rect 6229 6012 6293 6016
rect 6229 5956 6233 6012
rect 6233 5956 6289 6012
rect 6289 5956 6293 6012
rect 6229 5952 6293 5956
rect 6309 6012 6373 6016
rect 6309 5956 6313 6012
rect 6313 5956 6369 6012
rect 6369 5956 6373 6012
rect 6309 5952 6373 5956
rect 8116 6012 8180 6016
rect 8116 5956 8120 6012
rect 8120 5956 8176 6012
rect 8176 5956 8180 6012
rect 8116 5952 8180 5956
rect 8196 6012 8260 6016
rect 8196 5956 8200 6012
rect 8200 5956 8256 6012
rect 8256 5956 8260 6012
rect 8196 5952 8260 5956
rect 8276 6012 8340 6016
rect 8276 5956 8280 6012
rect 8280 5956 8336 6012
rect 8336 5956 8340 6012
rect 8276 5952 8340 5956
rect 8356 6012 8420 6016
rect 8356 5956 8360 6012
rect 8360 5956 8416 6012
rect 8416 5956 8420 6012
rect 8356 5952 8420 5956
rect 2635 5468 2699 5472
rect 2635 5412 2639 5468
rect 2639 5412 2695 5468
rect 2695 5412 2699 5468
rect 2635 5408 2699 5412
rect 2715 5468 2779 5472
rect 2715 5412 2719 5468
rect 2719 5412 2775 5468
rect 2775 5412 2779 5468
rect 2715 5408 2779 5412
rect 2795 5468 2859 5472
rect 2795 5412 2799 5468
rect 2799 5412 2855 5468
rect 2855 5412 2859 5468
rect 2795 5408 2859 5412
rect 2875 5468 2939 5472
rect 2875 5412 2879 5468
rect 2879 5412 2935 5468
rect 2935 5412 2939 5468
rect 2875 5408 2939 5412
rect 4682 5468 4746 5472
rect 4682 5412 4686 5468
rect 4686 5412 4742 5468
rect 4742 5412 4746 5468
rect 4682 5408 4746 5412
rect 4762 5468 4826 5472
rect 4762 5412 4766 5468
rect 4766 5412 4822 5468
rect 4822 5412 4826 5468
rect 4762 5408 4826 5412
rect 4842 5468 4906 5472
rect 4842 5412 4846 5468
rect 4846 5412 4902 5468
rect 4902 5412 4906 5468
rect 4842 5408 4906 5412
rect 4922 5468 4986 5472
rect 4922 5412 4926 5468
rect 4926 5412 4982 5468
rect 4982 5412 4986 5468
rect 4922 5408 4986 5412
rect 6729 5468 6793 5472
rect 6729 5412 6733 5468
rect 6733 5412 6789 5468
rect 6789 5412 6793 5468
rect 6729 5408 6793 5412
rect 6809 5468 6873 5472
rect 6809 5412 6813 5468
rect 6813 5412 6869 5468
rect 6869 5412 6873 5468
rect 6809 5408 6873 5412
rect 6889 5468 6953 5472
rect 6889 5412 6893 5468
rect 6893 5412 6949 5468
rect 6949 5412 6953 5468
rect 6889 5408 6953 5412
rect 6969 5468 7033 5472
rect 6969 5412 6973 5468
rect 6973 5412 7029 5468
rect 7029 5412 7033 5468
rect 6969 5408 7033 5412
rect 8776 5468 8840 5472
rect 8776 5412 8780 5468
rect 8780 5412 8836 5468
rect 8836 5412 8840 5468
rect 8776 5408 8840 5412
rect 8856 5468 8920 5472
rect 8856 5412 8860 5468
rect 8860 5412 8916 5468
rect 8916 5412 8920 5468
rect 8856 5408 8920 5412
rect 8936 5468 9000 5472
rect 8936 5412 8940 5468
rect 8940 5412 8996 5468
rect 8996 5412 9000 5468
rect 8936 5408 9000 5412
rect 9016 5468 9080 5472
rect 9016 5412 9020 5468
rect 9020 5412 9076 5468
rect 9076 5412 9080 5468
rect 9016 5408 9080 5412
rect 1975 4924 2039 4928
rect 1975 4868 1979 4924
rect 1979 4868 2035 4924
rect 2035 4868 2039 4924
rect 1975 4864 2039 4868
rect 2055 4924 2119 4928
rect 2055 4868 2059 4924
rect 2059 4868 2115 4924
rect 2115 4868 2119 4924
rect 2055 4864 2119 4868
rect 2135 4924 2199 4928
rect 2135 4868 2139 4924
rect 2139 4868 2195 4924
rect 2195 4868 2199 4924
rect 2135 4864 2199 4868
rect 2215 4924 2279 4928
rect 2215 4868 2219 4924
rect 2219 4868 2275 4924
rect 2275 4868 2279 4924
rect 2215 4864 2279 4868
rect 4022 4924 4086 4928
rect 4022 4868 4026 4924
rect 4026 4868 4082 4924
rect 4082 4868 4086 4924
rect 4022 4864 4086 4868
rect 4102 4924 4166 4928
rect 4102 4868 4106 4924
rect 4106 4868 4162 4924
rect 4162 4868 4166 4924
rect 4102 4864 4166 4868
rect 4182 4924 4246 4928
rect 4182 4868 4186 4924
rect 4186 4868 4242 4924
rect 4242 4868 4246 4924
rect 4182 4864 4246 4868
rect 4262 4924 4326 4928
rect 4262 4868 4266 4924
rect 4266 4868 4322 4924
rect 4322 4868 4326 4924
rect 4262 4864 4326 4868
rect 6069 4924 6133 4928
rect 6069 4868 6073 4924
rect 6073 4868 6129 4924
rect 6129 4868 6133 4924
rect 6069 4864 6133 4868
rect 6149 4924 6213 4928
rect 6149 4868 6153 4924
rect 6153 4868 6209 4924
rect 6209 4868 6213 4924
rect 6149 4864 6213 4868
rect 6229 4924 6293 4928
rect 6229 4868 6233 4924
rect 6233 4868 6289 4924
rect 6289 4868 6293 4924
rect 6229 4864 6293 4868
rect 6309 4924 6373 4928
rect 6309 4868 6313 4924
rect 6313 4868 6369 4924
rect 6369 4868 6373 4924
rect 6309 4864 6373 4868
rect 8116 4924 8180 4928
rect 8116 4868 8120 4924
rect 8120 4868 8176 4924
rect 8176 4868 8180 4924
rect 8116 4864 8180 4868
rect 8196 4924 8260 4928
rect 8196 4868 8200 4924
rect 8200 4868 8256 4924
rect 8256 4868 8260 4924
rect 8196 4864 8260 4868
rect 8276 4924 8340 4928
rect 8276 4868 8280 4924
rect 8280 4868 8336 4924
rect 8336 4868 8340 4924
rect 8276 4864 8340 4868
rect 8356 4924 8420 4928
rect 8356 4868 8360 4924
rect 8360 4868 8416 4924
rect 8416 4868 8420 4924
rect 8356 4864 8420 4868
rect 5764 4660 5828 4724
rect 2635 4380 2699 4384
rect 2635 4324 2639 4380
rect 2639 4324 2695 4380
rect 2695 4324 2699 4380
rect 2635 4320 2699 4324
rect 2715 4380 2779 4384
rect 2715 4324 2719 4380
rect 2719 4324 2775 4380
rect 2775 4324 2779 4380
rect 2715 4320 2779 4324
rect 2795 4380 2859 4384
rect 2795 4324 2799 4380
rect 2799 4324 2855 4380
rect 2855 4324 2859 4380
rect 2795 4320 2859 4324
rect 2875 4380 2939 4384
rect 2875 4324 2879 4380
rect 2879 4324 2935 4380
rect 2935 4324 2939 4380
rect 2875 4320 2939 4324
rect 4682 4380 4746 4384
rect 4682 4324 4686 4380
rect 4686 4324 4742 4380
rect 4742 4324 4746 4380
rect 4682 4320 4746 4324
rect 4762 4380 4826 4384
rect 4762 4324 4766 4380
rect 4766 4324 4822 4380
rect 4822 4324 4826 4380
rect 4762 4320 4826 4324
rect 4842 4380 4906 4384
rect 4842 4324 4846 4380
rect 4846 4324 4902 4380
rect 4902 4324 4906 4380
rect 4842 4320 4906 4324
rect 4922 4380 4986 4384
rect 4922 4324 4926 4380
rect 4926 4324 4982 4380
rect 4982 4324 4986 4380
rect 4922 4320 4986 4324
rect 6729 4380 6793 4384
rect 6729 4324 6733 4380
rect 6733 4324 6789 4380
rect 6789 4324 6793 4380
rect 6729 4320 6793 4324
rect 6809 4380 6873 4384
rect 6809 4324 6813 4380
rect 6813 4324 6869 4380
rect 6869 4324 6873 4380
rect 6809 4320 6873 4324
rect 6889 4380 6953 4384
rect 6889 4324 6893 4380
rect 6893 4324 6949 4380
rect 6949 4324 6953 4380
rect 6889 4320 6953 4324
rect 6969 4380 7033 4384
rect 6969 4324 6973 4380
rect 6973 4324 7029 4380
rect 7029 4324 7033 4380
rect 6969 4320 7033 4324
rect 8776 4380 8840 4384
rect 8776 4324 8780 4380
rect 8780 4324 8836 4380
rect 8836 4324 8840 4380
rect 8776 4320 8840 4324
rect 8856 4380 8920 4384
rect 8856 4324 8860 4380
rect 8860 4324 8916 4380
rect 8916 4324 8920 4380
rect 8856 4320 8920 4324
rect 8936 4380 9000 4384
rect 8936 4324 8940 4380
rect 8940 4324 8996 4380
rect 8996 4324 9000 4380
rect 8936 4320 9000 4324
rect 9016 4380 9080 4384
rect 9016 4324 9020 4380
rect 9020 4324 9076 4380
rect 9076 4324 9080 4380
rect 9016 4320 9080 4324
rect 1975 3836 2039 3840
rect 1975 3780 1979 3836
rect 1979 3780 2035 3836
rect 2035 3780 2039 3836
rect 1975 3776 2039 3780
rect 2055 3836 2119 3840
rect 2055 3780 2059 3836
rect 2059 3780 2115 3836
rect 2115 3780 2119 3836
rect 2055 3776 2119 3780
rect 2135 3836 2199 3840
rect 2135 3780 2139 3836
rect 2139 3780 2195 3836
rect 2195 3780 2199 3836
rect 2135 3776 2199 3780
rect 2215 3836 2279 3840
rect 2215 3780 2219 3836
rect 2219 3780 2275 3836
rect 2275 3780 2279 3836
rect 2215 3776 2279 3780
rect 4022 3836 4086 3840
rect 4022 3780 4026 3836
rect 4026 3780 4082 3836
rect 4082 3780 4086 3836
rect 4022 3776 4086 3780
rect 4102 3836 4166 3840
rect 4102 3780 4106 3836
rect 4106 3780 4162 3836
rect 4162 3780 4166 3836
rect 4102 3776 4166 3780
rect 4182 3836 4246 3840
rect 4182 3780 4186 3836
rect 4186 3780 4242 3836
rect 4242 3780 4246 3836
rect 4182 3776 4246 3780
rect 4262 3836 4326 3840
rect 4262 3780 4266 3836
rect 4266 3780 4322 3836
rect 4322 3780 4326 3836
rect 4262 3776 4326 3780
rect 6069 3836 6133 3840
rect 6069 3780 6073 3836
rect 6073 3780 6129 3836
rect 6129 3780 6133 3836
rect 6069 3776 6133 3780
rect 6149 3836 6213 3840
rect 6149 3780 6153 3836
rect 6153 3780 6209 3836
rect 6209 3780 6213 3836
rect 6149 3776 6213 3780
rect 6229 3836 6293 3840
rect 6229 3780 6233 3836
rect 6233 3780 6289 3836
rect 6289 3780 6293 3836
rect 6229 3776 6293 3780
rect 6309 3836 6373 3840
rect 6309 3780 6313 3836
rect 6313 3780 6369 3836
rect 6369 3780 6373 3836
rect 6309 3776 6373 3780
rect 8116 3836 8180 3840
rect 8116 3780 8120 3836
rect 8120 3780 8176 3836
rect 8176 3780 8180 3836
rect 8116 3776 8180 3780
rect 8196 3836 8260 3840
rect 8196 3780 8200 3836
rect 8200 3780 8256 3836
rect 8256 3780 8260 3836
rect 8196 3776 8260 3780
rect 8276 3836 8340 3840
rect 8276 3780 8280 3836
rect 8280 3780 8336 3836
rect 8336 3780 8340 3836
rect 8276 3776 8340 3780
rect 8356 3836 8420 3840
rect 8356 3780 8360 3836
rect 8360 3780 8416 3836
rect 8416 3780 8420 3836
rect 8356 3776 8420 3780
rect 2635 3292 2699 3296
rect 2635 3236 2639 3292
rect 2639 3236 2695 3292
rect 2695 3236 2699 3292
rect 2635 3232 2699 3236
rect 2715 3292 2779 3296
rect 2715 3236 2719 3292
rect 2719 3236 2775 3292
rect 2775 3236 2779 3292
rect 2715 3232 2779 3236
rect 2795 3292 2859 3296
rect 2795 3236 2799 3292
rect 2799 3236 2855 3292
rect 2855 3236 2859 3292
rect 2795 3232 2859 3236
rect 2875 3292 2939 3296
rect 2875 3236 2879 3292
rect 2879 3236 2935 3292
rect 2935 3236 2939 3292
rect 2875 3232 2939 3236
rect 4682 3292 4746 3296
rect 4682 3236 4686 3292
rect 4686 3236 4742 3292
rect 4742 3236 4746 3292
rect 4682 3232 4746 3236
rect 4762 3292 4826 3296
rect 4762 3236 4766 3292
rect 4766 3236 4822 3292
rect 4822 3236 4826 3292
rect 4762 3232 4826 3236
rect 4842 3292 4906 3296
rect 4842 3236 4846 3292
rect 4846 3236 4902 3292
rect 4902 3236 4906 3292
rect 4842 3232 4906 3236
rect 4922 3292 4986 3296
rect 4922 3236 4926 3292
rect 4926 3236 4982 3292
rect 4982 3236 4986 3292
rect 4922 3232 4986 3236
rect 6729 3292 6793 3296
rect 6729 3236 6733 3292
rect 6733 3236 6789 3292
rect 6789 3236 6793 3292
rect 6729 3232 6793 3236
rect 6809 3292 6873 3296
rect 6809 3236 6813 3292
rect 6813 3236 6869 3292
rect 6869 3236 6873 3292
rect 6809 3232 6873 3236
rect 6889 3292 6953 3296
rect 6889 3236 6893 3292
rect 6893 3236 6949 3292
rect 6949 3236 6953 3292
rect 6889 3232 6953 3236
rect 6969 3292 7033 3296
rect 6969 3236 6973 3292
rect 6973 3236 7029 3292
rect 7029 3236 7033 3292
rect 6969 3232 7033 3236
rect 8776 3292 8840 3296
rect 8776 3236 8780 3292
rect 8780 3236 8836 3292
rect 8836 3236 8840 3292
rect 8776 3232 8840 3236
rect 8856 3292 8920 3296
rect 8856 3236 8860 3292
rect 8860 3236 8916 3292
rect 8916 3236 8920 3292
rect 8856 3232 8920 3236
rect 8936 3292 9000 3296
rect 8936 3236 8940 3292
rect 8940 3236 8996 3292
rect 8996 3236 9000 3292
rect 8936 3232 9000 3236
rect 9016 3292 9080 3296
rect 9016 3236 9020 3292
rect 9020 3236 9076 3292
rect 9076 3236 9080 3292
rect 9016 3232 9080 3236
rect 1975 2748 2039 2752
rect 1975 2692 1979 2748
rect 1979 2692 2035 2748
rect 2035 2692 2039 2748
rect 1975 2688 2039 2692
rect 2055 2748 2119 2752
rect 2055 2692 2059 2748
rect 2059 2692 2115 2748
rect 2115 2692 2119 2748
rect 2055 2688 2119 2692
rect 2135 2748 2199 2752
rect 2135 2692 2139 2748
rect 2139 2692 2195 2748
rect 2195 2692 2199 2748
rect 2135 2688 2199 2692
rect 2215 2748 2279 2752
rect 2215 2692 2219 2748
rect 2219 2692 2275 2748
rect 2275 2692 2279 2748
rect 2215 2688 2279 2692
rect 4022 2748 4086 2752
rect 4022 2692 4026 2748
rect 4026 2692 4082 2748
rect 4082 2692 4086 2748
rect 4022 2688 4086 2692
rect 4102 2748 4166 2752
rect 4102 2692 4106 2748
rect 4106 2692 4162 2748
rect 4162 2692 4166 2748
rect 4102 2688 4166 2692
rect 4182 2748 4246 2752
rect 4182 2692 4186 2748
rect 4186 2692 4242 2748
rect 4242 2692 4246 2748
rect 4182 2688 4246 2692
rect 4262 2748 4326 2752
rect 4262 2692 4266 2748
rect 4266 2692 4322 2748
rect 4322 2692 4326 2748
rect 4262 2688 4326 2692
rect 6069 2748 6133 2752
rect 6069 2692 6073 2748
rect 6073 2692 6129 2748
rect 6129 2692 6133 2748
rect 6069 2688 6133 2692
rect 6149 2748 6213 2752
rect 6149 2692 6153 2748
rect 6153 2692 6209 2748
rect 6209 2692 6213 2748
rect 6149 2688 6213 2692
rect 6229 2748 6293 2752
rect 6229 2692 6233 2748
rect 6233 2692 6289 2748
rect 6289 2692 6293 2748
rect 6229 2688 6293 2692
rect 6309 2748 6373 2752
rect 6309 2692 6313 2748
rect 6313 2692 6369 2748
rect 6369 2692 6373 2748
rect 6309 2688 6373 2692
rect 8116 2748 8180 2752
rect 8116 2692 8120 2748
rect 8120 2692 8176 2748
rect 8176 2692 8180 2748
rect 8116 2688 8180 2692
rect 8196 2748 8260 2752
rect 8196 2692 8200 2748
rect 8200 2692 8256 2748
rect 8256 2692 8260 2748
rect 8196 2688 8260 2692
rect 8276 2748 8340 2752
rect 8276 2692 8280 2748
rect 8280 2692 8336 2748
rect 8336 2692 8340 2748
rect 8276 2688 8340 2692
rect 8356 2748 8420 2752
rect 8356 2692 8360 2748
rect 8360 2692 8416 2748
rect 8416 2692 8420 2748
rect 8356 2688 8420 2692
rect 2635 2204 2699 2208
rect 2635 2148 2639 2204
rect 2639 2148 2695 2204
rect 2695 2148 2699 2204
rect 2635 2144 2699 2148
rect 2715 2204 2779 2208
rect 2715 2148 2719 2204
rect 2719 2148 2775 2204
rect 2775 2148 2779 2204
rect 2715 2144 2779 2148
rect 2795 2204 2859 2208
rect 2795 2148 2799 2204
rect 2799 2148 2855 2204
rect 2855 2148 2859 2204
rect 2795 2144 2859 2148
rect 2875 2204 2939 2208
rect 2875 2148 2879 2204
rect 2879 2148 2935 2204
rect 2935 2148 2939 2204
rect 2875 2144 2939 2148
rect 4682 2204 4746 2208
rect 4682 2148 4686 2204
rect 4686 2148 4742 2204
rect 4742 2148 4746 2204
rect 4682 2144 4746 2148
rect 4762 2204 4826 2208
rect 4762 2148 4766 2204
rect 4766 2148 4822 2204
rect 4822 2148 4826 2204
rect 4762 2144 4826 2148
rect 4842 2204 4906 2208
rect 4842 2148 4846 2204
rect 4846 2148 4902 2204
rect 4902 2148 4906 2204
rect 4842 2144 4906 2148
rect 4922 2204 4986 2208
rect 4922 2148 4926 2204
rect 4926 2148 4982 2204
rect 4982 2148 4986 2204
rect 4922 2144 4986 2148
rect 6729 2204 6793 2208
rect 6729 2148 6733 2204
rect 6733 2148 6789 2204
rect 6789 2148 6793 2204
rect 6729 2144 6793 2148
rect 6809 2204 6873 2208
rect 6809 2148 6813 2204
rect 6813 2148 6869 2204
rect 6869 2148 6873 2204
rect 6809 2144 6873 2148
rect 6889 2204 6953 2208
rect 6889 2148 6893 2204
rect 6893 2148 6949 2204
rect 6949 2148 6953 2204
rect 6889 2144 6953 2148
rect 6969 2204 7033 2208
rect 6969 2148 6973 2204
rect 6973 2148 7029 2204
rect 7029 2148 7033 2204
rect 6969 2144 7033 2148
rect 8776 2204 8840 2208
rect 8776 2148 8780 2204
rect 8780 2148 8836 2204
rect 8836 2148 8840 2204
rect 8776 2144 8840 2148
rect 8856 2204 8920 2208
rect 8856 2148 8860 2204
rect 8860 2148 8916 2204
rect 8916 2148 8920 2204
rect 8856 2144 8920 2148
rect 8936 2204 9000 2208
rect 8936 2148 8940 2204
rect 8940 2148 8996 2204
rect 8996 2148 9000 2204
rect 8936 2144 9000 2148
rect 9016 2204 9080 2208
rect 9016 2148 9020 2204
rect 9020 2148 9076 2204
rect 9076 2148 9080 2204
rect 9016 2144 9080 2148
<< metal4 >>
rect 1967 10368 2287 10384
rect 1967 10304 1975 10368
rect 2039 10304 2055 10368
rect 2119 10304 2135 10368
rect 2199 10304 2215 10368
rect 2279 10304 2287 10368
rect 1967 9434 2287 10304
rect 1967 9280 2009 9434
rect 2245 9280 2287 9434
rect 1967 9216 1975 9280
rect 2279 9216 2287 9280
rect 1967 9198 2009 9216
rect 2245 9198 2287 9216
rect 1967 8192 2287 9198
rect 1967 8128 1975 8192
rect 2039 8128 2055 8192
rect 2119 8128 2135 8192
rect 2199 8128 2215 8192
rect 2279 8128 2287 8192
rect 1967 7394 2287 8128
rect 1967 7158 2009 7394
rect 2245 7158 2287 7394
rect 1967 7104 2287 7158
rect 1967 7040 1975 7104
rect 2039 7040 2055 7104
rect 2119 7040 2135 7104
rect 2199 7040 2215 7104
rect 2279 7040 2287 7104
rect 1967 6016 2287 7040
rect 1967 5952 1975 6016
rect 2039 5952 2055 6016
rect 2119 5952 2135 6016
rect 2199 5952 2215 6016
rect 2279 5952 2287 6016
rect 1967 5354 2287 5952
rect 1967 5118 2009 5354
rect 2245 5118 2287 5354
rect 1967 4928 2287 5118
rect 1967 4864 1975 4928
rect 2039 4864 2055 4928
rect 2119 4864 2135 4928
rect 2199 4864 2215 4928
rect 2279 4864 2287 4928
rect 1967 3840 2287 4864
rect 1967 3776 1975 3840
rect 2039 3776 2055 3840
rect 2119 3776 2135 3840
rect 2199 3776 2215 3840
rect 2279 3776 2287 3840
rect 1967 3314 2287 3776
rect 1967 3078 2009 3314
rect 2245 3078 2287 3314
rect 1967 2752 2287 3078
rect 1967 2688 1975 2752
rect 2039 2688 2055 2752
rect 2119 2688 2135 2752
rect 2199 2688 2215 2752
rect 2279 2688 2287 2752
rect 1967 2128 2287 2688
rect 2627 10094 2947 10384
rect 2627 9858 2669 10094
rect 2905 9858 2947 10094
rect 2627 9824 2947 9858
rect 2627 9760 2635 9824
rect 2699 9760 2715 9824
rect 2779 9760 2795 9824
rect 2859 9760 2875 9824
rect 2939 9760 2947 9824
rect 2627 8736 2947 9760
rect 2627 8672 2635 8736
rect 2699 8672 2715 8736
rect 2779 8672 2795 8736
rect 2859 8672 2875 8736
rect 2939 8672 2947 8736
rect 2627 8054 2947 8672
rect 2627 7818 2669 8054
rect 2905 7818 2947 8054
rect 2627 7648 2947 7818
rect 2627 7584 2635 7648
rect 2699 7584 2715 7648
rect 2779 7584 2795 7648
rect 2859 7584 2875 7648
rect 2939 7584 2947 7648
rect 2627 6560 2947 7584
rect 2627 6496 2635 6560
rect 2699 6496 2715 6560
rect 2779 6496 2795 6560
rect 2859 6496 2875 6560
rect 2939 6496 2947 6560
rect 2627 6014 2947 6496
rect 2627 5778 2669 6014
rect 2905 5778 2947 6014
rect 2627 5472 2947 5778
rect 2627 5408 2635 5472
rect 2699 5408 2715 5472
rect 2779 5408 2795 5472
rect 2859 5408 2875 5472
rect 2939 5408 2947 5472
rect 2627 4384 2947 5408
rect 2627 4320 2635 4384
rect 2699 4320 2715 4384
rect 2779 4320 2795 4384
rect 2859 4320 2875 4384
rect 2939 4320 2947 4384
rect 2627 3974 2947 4320
rect 2627 3738 2669 3974
rect 2905 3738 2947 3974
rect 2627 3296 2947 3738
rect 2627 3232 2635 3296
rect 2699 3232 2715 3296
rect 2779 3232 2795 3296
rect 2859 3232 2875 3296
rect 2939 3232 2947 3296
rect 2627 2208 2947 3232
rect 2627 2144 2635 2208
rect 2699 2144 2715 2208
rect 2779 2144 2795 2208
rect 2859 2144 2875 2208
rect 2939 2144 2947 2208
rect 2627 2128 2947 2144
rect 4014 10368 4334 10384
rect 4014 10304 4022 10368
rect 4086 10304 4102 10368
rect 4166 10304 4182 10368
rect 4246 10304 4262 10368
rect 4326 10304 4334 10368
rect 4014 9434 4334 10304
rect 4014 9280 4056 9434
rect 4292 9280 4334 9434
rect 4014 9216 4022 9280
rect 4326 9216 4334 9280
rect 4014 9198 4056 9216
rect 4292 9198 4334 9216
rect 4014 8192 4334 9198
rect 4014 8128 4022 8192
rect 4086 8128 4102 8192
rect 4166 8128 4182 8192
rect 4246 8128 4262 8192
rect 4326 8128 4334 8192
rect 4014 7394 4334 8128
rect 4014 7158 4056 7394
rect 4292 7158 4334 7394
rect 4014 7104 4334 7158
rect 4014 7040 4022 7104
rect 4086 7040 4102 7104
rect 4166 7040 4182 7104
rect 4246 7040 4262 7104
rect 4326 7040 4334 7104
rect 4014 6016 4334 7040
rect 4014 5952 4022 6016
rect 4086 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4334 6016
rect 4014 5354 4334 5952
rect 4014 5118 4056 5354
rect 4292 5118 4334 5354
rect 4014 4928 4334 5118
rect 4014 4864 4022 4928
rect 4086 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4334 4928
rect 4014 3840 4334 4864
rect 4014 3776 4022 3840
rect 4086 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4334 3840
rect 4014 3314 4334 3776
rect 4014 3078 4056 3314
rect 4292 3078 4334 3314
rect 4014 2752 4334 3078
rect 4014 2688 4022 2752
rect 4086 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4334 2752
rect 4014 2128 4334 2688
rect 4674 10094 4994 10384
rect 4674 9858 4716 10094
rect 4952 9858 4994 10094
rect 4674 9824 4994 9858
rect 4674 9760 4682 9824
rect 4746 9760 4762 9824
rect 4826 9760 4842 9824
rect 4906 9760 4922 9824
rect 4986 9760 4994 9824
rect 4674 8736 4994 9760
rect 4674 8672 4682 8736
rect 4746 8672 4762 8736
rect 4826 8672 4842 8736
rect 4906 8672 4922 8736
rect 4986 8672 4994 8736
rect 4674 8054 4994 8672
rect 4674 7818 4716 8054
rect 4952 7818 4994 8054
rect 4674 7648 4994 7818
rect 4674 7584 4682 7648
rect 4746 7584 4762 7648
rect 4826 7584 4842 7648
rect 4906 7584 4922 7648
rect 4986 7584 4994 7648
rect 4674 6560 4994 7584
rect 6061 10368 6381 10384
rect 6061 10304 6069 10368
rect 6133 10304 6149 10368
rect 6213 10304 6229 10368
rect 6293 10304 6309 10368
rect 6373 10304 6381 10368
rect 6061 9434 6381 10304
rect 6061 9280 6103 9434
rect 6339 9280 6381 9434
rect 6061 9216 6069 9280
rect 6373 9216 6381 9280
rect 6061 9198 6103 9216
rect 6339 9198 6381 9216
rect 6061 8192 6381 9198
rect 6061 8128 6069 8192
rect 6133 8128 6149 8192
rect 6213 8128 6229 8192
rect 6293 8128 6309 8192
rect 6373 8128 6381 8192
rect 5763 7444 5829 7445
rect 5763 7380 5764 7444
rect 5828 7380 5829 7444
rect 5763 7379 5829 7380
rect 6061 7394 6381 8128
rect 4674 6496 4682 6560
rect 4746 6496 4762 6560
rect 4826 6496 4842 6560
rect 4906 6496 4922 6560
rect 4986 6496 4994 6560
rect 4674 6014 4994 6496
rect 4674 5778 4716 6014
rect 4952 5778 4994 6014
rect 4674 5472 4994 5778
rect 4674 5408 4682 5472
rect 4746 5408 4762 5472
rect 4826 5408 4842 5472
rect 4906 5408 4922 5472
rect 4986 5408 4994 5472
rect 4674 4384 4994 5408
rect 5766 4725 5826 7379
rect 6061 7158 6103 7394
rect 6339 7158 6381 7394
rect 6061 7104 6381 7158
rect 6061 7040 6069 7104
rect 6133 7040 6149 7104
rect 6213 7040 6229 7104
rect 6293 7040 6309 7104
rect 6373 7040 6381 7104
rect 6061 6016 6381 7040
rect 6061 5952 6069 6016
rect 6133 5952 6149 6016
rect 6213 5952 6229 6016
rect 6293 5952 6309 6016
rect 6373 5952 6381 6016
rect 6061 5354 6381 5952
rect 6061 5118 6103 5354
rect 6339 5118 6381 5354
rect 6061 4928 6381 5118
rect 6061 4864 6069 4928
rect 6133 4864 6149 4928
rect 6213 4864 6229 4928
rect 6293 4864 6309 4928
rect 6373 4864 6381 4928
rect 5763 4724 5829 4725
rect 5763 4660 5764 4724
rect 5828 4660 5829 4724
rect 5763 4659 5829 4660
rect 4674 4320 4682 4384
rect 4746 4320 4762 4384
rect 4826 4320 4842 4384
rect 4906 4320 4922 4384
rect 4986 4320 4994 4384
rect 4674 3974 4994 4320
rect 4674 3738 4716 3974
rect 4952 3738 4994 3974
rect 4674 3296 4994 3738
rect 4674 3232 4682 3296
rect 4746 3232 4762 3296
rect 4826 3232 4842 3296
rect 4906 3232 4922 3296
rect 4986 3232 4994 3296
rect 4674 2208 4994 3232
rect 4674 2144 4682 2208
rect 4746 2144 4762 2208
rect 4826 2144 4842 2208
rect 4906 2144 4922 2208
rect 4986 2144 4994 2208
rect 4674 2128 4994 2144
rect 6061 3840 6381 4864
rect 6061 3776 6069 3840
rect 6133 3776 6149 3840
rect 6213 3776 6229 3840
rect 6293 3776 6309 3840
rect 6373 3776 6381 3840
rect 6061 3314 6381 3776
rect 6061 3078 6103 3314
rect 6339 3078 6381 3314
rect 6061 2752 6381 3078
rect 6061 2688 6069 2752
rect 6133 2688 6149 2752
rect 6213 2688 6229 2752
rect 6293 2688 6309 2752
rect 6373 2688 6381 2752
rect 6061 2128 6381 2688
rect 6721 10094 7041 10384
rect 6721 9858 6763 10094
rect 6999 9858 7041 10094
rect 6721 9824 7041 9858
rect 6721 9760 6729 9824
rect 6793 9760 6809 9824
rect 6873 9760 6889 9824
rect 6953 9760 6969 9824
rect 7033 9760 7041 9824
rect 6721 8736 7041 9760
rect 6721 8672 6729 8736
rect 6793 8672 6809 8736
rect 6873 8672 6889 8736
rect 6953 8672 6969 8736
rect 7033 8672 7041 8736
rect 6721 8054 7041 8672
rect 6721 7818 6763 8054
rect 6999 7818 7041 8054
rect 6721 7648 7041 7818
rect 6721 7584 6729 7648
rect 6793 7584 6809 7648
rect 6873 7584 6889 7648
rect 6953 7584 6969 7648
rect 7033 7584 7041 7648
rect 6721 6560 7041 7584
rect 6721 6496 6729 6560
rect 6793 6496 6809 6560
rect 6873 6496 6889 6560
rect 6953 6496 6969 6560
rect 7033 6496 7041 6560
rect 6721 6014 7041 6496
rect 6721 5778 6763 6014
rect 6999 5778 7041 6014
rect 6721 5472 7041 5778
rect 6721 5408 6729 5472
rect 6793 5408 6809 5472
rect 6873 5408 6889 5472
rect 6953 5408 6969 5472
rect 7033 5408 7041 5472
rect 6721 4384 7041 5408
rect 6721 4320 6729 4384
rect 6793 4320 6809 4384
rect 6873 4320 6889 4384
rect 6953 4320 6969 4384
rect 7033 4320 7041 4384
rect 6721 3974 7041 4320
rect 6721 3738 6763 3974
rect 6999 3738 7041 3974
rect 6721 3296 7041 3738
rect 6721 3232 6729 3296
rect 6793 3232 6809 3296
rect 6873 3232 6889 3296
rect 6953 3232 6969 3296
rect 7033 3232 7041 3296
rect 6721 2208 7041 3232
rect 6721 2144 6729 2208
rect 6793 2144 6809 2208
rect 6873 2144 6889 2208
rect 6953 2144 6969 2208
rect 7033 2144 7041 2208
rect 6721 2128 7041 2144
rect 8108 10368 8428 10384
rect 8108 10304 8116 10368
rect 8180 10304 8196 10368
rect 8260 10304 8276 10368
rect 8340 10304 8356 10368
rect 8420 10304 8428 10368
rect 8108 9434 8428 10304
rect 8108 9280 8150 9434
rect 8386 9280 8428 9434
rect 8108 9216 8116 9280
rect 8420 9216 8428 9280
rect 8108 9198 8150 9216
rect 8386 9198 8428 9216
rect 8108 8192 8428 9198
rect 8108 8128 8116 8192
rect 8180 8128 8196 8192
rect 8260 8128 8276 8192
rect 8340 8128 8356 8192
rect 8420 8128 8428 8192
rect 8108 7394 8428 8128
rect 8108 7158 8150 7394
rect 8386 7158 8428 7394
rect 8108 7104 8428 7158
rect 8108 7040 8116 7104
rect 8180 7040 8196 7104
rect 8260 7040 8276 7104
rect 8340 7040 8356 7104
rect 8420 7040 8428 7104
rect 8108 6016 8428 7040
rect 8108 5952 8116 6016
rect 8180 5952 8196 6016
rect 8260 5952 8276 6016
rect 8340 5952 8356 6016
rect 8420 5952 8428 6016
rect 8108 5354 8428 5952
rect 8108 5118 8150 5354
rect 8386 5118 8428 5354
rect 8108 4928 8428 5118
rect 8108 4864 8116 4928
rect 8180 4864 8196 4928
rect 8260 4864 8276 4928
rect 8340 4864 8356 4928
rect 8420 4864 8428 4928
rect 8108 3840 8428 4864
rect 8108 3776 8116 3840
rect 8180 3776 8196 3840
rect 8260 3776 8276 3840
rect 8340 3776 8356 3840
rect 8420 3776 8428 3840
rect 8108 3314 8428 3776
rect 8108 3078 8150 3314
rect 8386 3078 8428 3314
rect 8108 2752 8428 3078
rect 8108 2688 8116 2752
rect 8180 2688 8196 2752
rect 8260 2688 8276 2752
rect 8340 2688 8356 2752
rect 8420 2688 8428 2752
rect 8108 2128 8428 2688
rect 8768 10094 9088 10384
rect 8768 9858 8810 10094
rect 9046 9858 9088 10094
rect 8768 9824 9088 9858
rect 8768 9760 8776 9824
rect 8840 9760 8856 9824
rect 8920 9760 8936 9824
rect 9000 9760 9016 9824
rect 9080 9760 9088 9824
rect 8768 8736 9088 9760
rect 8768 8672 8776 8736
rect 8840 8672 8856 8736
rect 8920 8672 8936 8736
rect 9000 8672 9016 8736
rect 9080 8672 9088 8736
rect 8768 8054 9088 8672
rect 8768 7818 8810 8054
rect 9046 7818 9088 8054
rect 8768 7648 9088 7818
rect 8768 7584 8776 7648
rect 8840 7584 8856 7648
rect 8920 7584 8936 7648
rect 9000 7584 9016 7648
rect 9080 7584 9088 7648
rect 8768 6560 9088 7584
rect 8768 6496 8776 6560
rect 8840 6496 8856 6560
rect 8920 6496 8936 6560
rect 9000 6496 9016 6560
rect 9080 6496 9088 6560
rect 8768 6014 9088 6496
rect 8768 5778 8810 6014
rect 9046 5778 9088 6014
rect 8768 5472 9088 5778
rect 8768 5408 8776 5472
rect 8840 5408 8856 5472
rect 8920 5408 8936 5472
rect 9000 5408 9016 5472
rect 9080 5408 9088 5472
rect 8768 4384 9088 5408
rect 8768 4320 8776 4384
rect 8840 4320 8856 4384
rect 8920 4320 8936 4384
rect 9000 4320 9016 4384
rect 9080 4320 9088 4384
rect 8768 3974 9088 4320
rect 8768 3738 8810 3974
rect 9046 3738 9088 3974
rect 8768 3296 9088 3738
rect 8768 3232 8776 3296
rect 8840 3232 8856 3296
rect 8920 3232 8936 3296
rect 9000 3232 9016 3296
rect 9080 3232 9088 3296
rect 8768 2208 9088 3232
rect 8768 2144 8776 2208
rect 8840 2144 8856 2208
rect 8920 2144 8936 2208
rect 9000 2144 9016 2208
rect 9080 2144 9088 2208
rect 8768 2128 9088 2144
<< via4 >>
rect 2009 9280 2245 9434
rect 2009 9216 2039 9280
rect 2039 9216 2055 9280
rect 2055 9216 2119 9280
rect 2119 9216 2135 9280
rect 2135 9216 2199 9280
rect 2199 9216 2215 9280
rect 2215 9216 2245 9280
rect 2009 9198 2245 9216
rect 2009 7158 2245 7394
rect 2009 5118 2245 5354
rect 2009 3078 2245 3314
rect 2669 9858 2905 10094
rect 2669 7818 2905 8054
rect 2669 5778 2905 6014
rect 2669 3738 2905 3974
rect 4056 9280 4292 9434
rect 4056 9216 4086 9280
rect 4086 9216 4102 9280
rect 4102 9216 4166 9280
rect 4166 9216 4182 9280
rect 4182 9216 4246 9280
rect 4246 9216 4262 9280
rect 4262 9216 4292 9280
rect 4056 9198 4292 9216
rect 4056 7158 4292 7394
rect 4056 5118 4292 5354
rect 4056 3078 4292 3314
rect 4716 9858 4952 10094
rect 4716 7818 4952 8054
rect 6103 9280 6339 9434
rect 6103 9216 6133 9280
rect 6133 9216 6149 9280
rect 6149 9216 6213 9280
rect 6213 9216 6229 9280
rect 6229 9216 6293 9280
rect 6293 9216 6309 9280
rect 6309 9216 6339 9280
rect 6103 9198 6339 9216
rect 4716 5778 4952 6014
rect 6103 7158 6339 7394
rect 6103 5118 6339 5354
rect 4716 3738 4952 3974
rect 6103 3078 6339 3314
rect 6763 9858 6999 10094
rect 6763 7818 6999 8054
rect 6763 5778 6999 6014
rect 6763 3738 6999 3974
rect 8150 9280 8386 9434
rect 8150 9216 8180 9280
rect 8180 9216 8196 9280
rect 8196 9216 8260 9280
rect 8260 9216 8276 9280
rect 8276 9216 8340 9280
rect 8340 9216 8356 9280
rect 8356 9216 8386 9280
rect 8150 9198 8386 9216
rect 8150 7158 8386 7394
rect 8150 5118 8386 5354
rect 8150 3078 8386 3314
rect 8810 9858 9046 10094
rect 8810 7818 9046 8054
rect 8810 5778 9046 6014
rect 8810 3738 9046 3974
<< metal5 >>
rect 1056 10094 9340 10136
rect 1056 9858 2669 10094
rect 2905 9858 4716 10094
rect 4952 9858 6763 10094
rect 6999 9858 8810 10094
rect 9046 9858 9340 10094
rect 1056 9816 9340 9858
rect 1056 9434 9340 9476
rect 1056 9198 2009 9434
rect 2245 9198 4056 9434
rect 4292 9198 6103 9434
rect 6339 9198 8150 9434
rect 8386 9198 9340 9434
rect 1056 9156 9340 9198
rect 1056 8054 9340 8096
rect 1056 7818 2669 8054
rect 2905 7818 4716 8054
rect 4952 7818 6763 8054
rect 6999 7818 8810 8054
rect 9046 7818 9340 8054
rect 1056 7776 9340 7818
rect 1056 7394 9340 7436
rect 1056 7158 2009 7394
rect 2245 7158 4056 7394
rect 4292 7158 6103 7394
rect 6339 7158 8150 7394
rect 8386 7158 9340 7394
rect 1056 7116 9340 7158
rect 1056 6014 9340 6056
rect 1056 5778 2669 6014
rect 2905 5778 4716 6014
rect 4952 5778 6763 6014
rect 6999 5778 8810 6014
rect 9046 5778 9340 6014
rect 1056 5736 9340 5778
rect 1056 5354 9340 5396
rect 1056 5118 2009 5354
rect 2245 5118 4056 5354
rect 4292 5118 6103 5354
rect 6339 5118 8150 5354
rect 8386 5118 9340 5354
rect 1056 5076 9340 5118
rect 1056 3974 9340 4016
rect 1056 3738 2669 3974
rect 2905 3738 4716 3974
rect 4952 3738 6763 3974
rect 6999 3738 8810 3974
rect 9046 3738 9340 3974
rect 1056 3696 9340 3738
rect 1056 3314 9340 3356
rect 1056 3078 2009 3314
rect 2245 3078 4056 3314
rect 4292 3078 6103 3314
rect 6339 3078 8150 3314
rect 8386 3078 9340 3314
rect 1056 3036 9340 3078
use sky130_fd_sc_hd__nand2_1  _103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6256 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _104_
timestamp 1694700623
transform -1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 4048 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _106_
timestamp 1694700623
transform -1 0 3680 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_4  _107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2852 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_2  _108_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _109_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 4692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _110_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3956 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _111_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6348 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__o2111ai_2  _112_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6808 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_2  _114_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6348 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _115_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 8280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _116_
timestamp 1694700623
transform -1 0 8280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _117_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 7176 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _118_
timestamp 1694700623
transform 1 0 2852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _120_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 8188 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _121_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6164 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2ai_1  _122_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 6256 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _123_
timestamp 1694700623
transform -1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_1  _124_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5336 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand4b_2  _125_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__nand3_1  _126_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _127_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _128_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 8188 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand4b_1  _129_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6348 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _130_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _131_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 8188 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _132_
timestamp 1694700623
transform 1 0 7912 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand4b_1  _133_
timestamp 1694700623
transform -1 0 7544 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2ai_1  _134_
timestamp 1694700623
transform -1 0 6900 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _135_
timestamp 1694700623
transform 1 0 7084 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _136_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 5520 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _137_
timestamp 1694700623
transform -1 0 5520 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_2  _138_
timestamp 1694700623
transform 1 0 5612 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _139_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2392 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_2  _140_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3036 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_2  _141_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4140 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__a32oi_4  _142_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4232 0 -1 5440
box -38 -48 2062 592
use sky130_fd_sc_hd__o21ai_1  _143_
timestamp 1694700623
transform 1 0 6716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _144_
timestamp 1694700623
transform 1 0 5704 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a32oi_1  _145_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 5704 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _146_
timestamp 1694700623
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 2668 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _148_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _149_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6348 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _150_
timestamp 1694700623
transform 1 0 2944 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _151_
timestamp 1694700623
transform -1 0 1932 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _152_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1380 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _153_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2760 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _154_
timestamp 1694700623
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _155_
timestamp 1694700623
transform 1 0 3496 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _156_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1748 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_1  _157_
timestamp 1694700623
transform 1 0 1380 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _158_
timestamp 1694700623
transform 1 0 2944 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _159_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _160_
timestamp 1694700623
transform 1 0 4508 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _161_
timestamp 1694700623
transform 1 0 2852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _162_
timestamp 1694700623
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _163_
timestamp 1694700623
transform 1 0 1564 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3036 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _165_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4692 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _166_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _167_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 4416 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1694700623
transform -1 0 8280 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _169_
timestamp 1694700623
transform 1 0 7360 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _170_
timestamp 1694700623
transform -1 0 7268 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _171_
timestamp 1694700623
transform 1 0 7268 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _172_
timestamp 1694700623
transform 1 0 6440 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6808 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _174_
timestamp 1694700623
transform 1 0 7636 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _175_
timestamp 1694700623
transform -1 0 6900 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _176_
timestamp 1694700623
transform -1 0 8096 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1694700623
transform -1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 7728 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2ai_1  _179_
timestamp 1694700623
transform 1 0 6900 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp 1694700623
transform -1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_2  _181_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3772 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _182_
timestamp 1694700623
transform -1 0 4140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_1  _183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5060 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _184_
timestamp 1694700623
transform -1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1694700623
transform -1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _186_
timestamp 1694700623
transform -1 0 2760 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _187_
timestamp 1694700623
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _188_
timestamp 1694700623
transform 1 0 3864 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  _189_
timestamp 1694700623
transform -1 0 4508 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _190_
timestamp 1694700623
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_2  _191_
timestamp 1694700623
transform 1 0 5152 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _192_
timestamp 1694700623
transform -1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _193_
timestamp 1694700623
transform 1 0 4048 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__o2111ai_1  _194_
timestamp 1694700623
transform -1 0 5152 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2ai_1  _195_
timestamp 1694700623
transform 1 0 5336 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4692 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _197_
timestamp 1694700623
transform 1 0 4508 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _198_
timestamp 1694700623
transform -1 0 2852 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_4  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3588 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _200_
timestamp 1694700623
transform 1 0 7268 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _201_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5704 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _202_
timestamp 1694700623
transform 1 0 8556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _203_
timestamp 1694700623
transform -1 0 2392 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _204_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 7728 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _205_
timestamp 1694700623
transform -1 0 6716 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _206_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7452 0 -1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _207_
timestamp 1694700623
transform 1 0 6348 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _208_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 7360 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _209_
timestamp 1694700623
transform 1 0 6624 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _210_
timestamp 1694700623
transform 1 0 4784 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _211_
timestamp 1694700623
transform 1 0 1380 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _212_
timestamp 1694700623
transform 1 0 1380 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _213_
timestamp 1694700623
transform 1 0 1380 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _214_
timestamp 1694700623
transform 1 0 1380 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _215_
timestamp 1694700623
transform 1 0 1840 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _216_
timestamp 1694700623
transform 1 0 3312 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _217_
timestamp 1694700623
transform 1 0 7360 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _218_
timestamp 1694700623
transform 1 0 7544 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _219_
timestamp 1694700623
transform 1 0 1380 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _220_
timestamp 1694700623
transform 1 0 1564 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _221_
timestamp 1694700623
transform -1 0 6072 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4416 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1694700623
transform -1 0 5520 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1694700623
transform 1 0 4416 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clone2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_19
timestamp 1694700623
transform 1 0 2852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37
timestamp 1694700623
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_76 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 8096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1694700623
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_3
timestamp 1694700623
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_37
timestamp 1694700623
transform 1 0 4508 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1694700623
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_82 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_7
timestamp 1694700623
transform 1 0 1748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_26
timestamp 1694700623
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_29
timestamp 1694700623
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_54
timestamp 1694700623
transform 1 0 6072 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_63
timestamp 1694700623
transform 1 0 6900 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_81
timestamp 1694700623
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_85
timestamp 1694700623
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_27
timestamp 1694700623
transform 1 0 3588 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_48
timestamp 1694700623
transform 1 0 5520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 1694700623
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_72
timestamp 1694700623
transform 1 0 7728 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_81
timestamp 1694700623
transform 1 0 8556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_85
timestamp 1694700623
transform 1 0 8924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_3
timestamp 1694700623
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_29
timestamp 1694700623
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_61
timestamp 1694700623
transform 1 0 6716 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 1694700623
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_85
timestamp 1694700623
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_32
timestamp 1694700623
transform 1 0 4048 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_71
timestamp 1694700623
transform 1 0 7636 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_84
timestamp 1694700623
transform 1 0 8832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_29
timestamp 1694700623
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_55
timestamp 1694700623
transform 1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1694700623
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_85
timestamp 1694700623
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_17
timestamp 1694700623
transform 1 0 2668 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_64
timestamp 1694700623
transform 1 0 6992 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_39
timestamp 1694700623
transform 1 0 4692 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_85
timestamp 1694700623
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_44
timestamp 1694700623
transform 1 0 5152 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_85
timestamp 1694700623
transform 1 0 8924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 1694700623
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_18
timestamp 1694700623
transform 1 0 2760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 4048 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_38
timestamp 1694700623
transform 1 0 4600 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_47
timestamp 1694700623
transform 1 0 5428 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_79
timestamp 1694700623
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1694700623
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_85
timestamp 1694700623
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_27
timestamp 1694700623
transform 1 0 3588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1694700623
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_42
timestamp 1694700623
transform 1 0 4968 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_55
timestamp 1694700623
transform 1 0 6164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_72
timestamp 1694700623
transform 1 0 7728 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1694700623
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 1694700623
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_84
timestamp 1694700623
transform 1 0 8832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_3
timestamp 1694700623
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_11
timestamp 1694700623
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_19
timestamp 1694700623
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1694700623
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_40
timestamp 1694700623
transform 1 0 4784 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_48
timestamp 1694700623
transform 1 0 5520 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_63
timestamp 1694700623
transform 1 0 6900 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_78
timestamp 1694700623
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 1694700623
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform -1 0 7084 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1694700623
transform 1 0 4600 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1694700623
transform -1 0 3496 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1694700623
transform -1 0 8740 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1694700623
transform -1 0 4508 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1694700623
transform -1 0 3588 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1694700623
transform -1 0 8648 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1694700623
transform -1 0 7728 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1694700623
transform -1 0 8924 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1694700623
transform -1 0 2852 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1694700623
transform -1 0 8188 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1694700623
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1694700623
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output4
timestamp 1694700623
transform -1 0 6900 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_15
timestamp 1694700623
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1694700623
transform -1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_16
timestamp 1694700623
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1694700623
transform -1 0 9292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_17
timestamp 1694700623
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1694700623
transform -1 0 9292 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_18
timestamp 1694700623
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1694700623
transform -1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_19
timestamp 1694700623
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1694700623
transform -1 0 9292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_20
timestamp 1694700623
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1694700623
transform -1 0 9292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_21
timestamp 1694700623
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1694700623
transform -1 0 9292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_22
timestamp 1694700623
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1694700623
transform -1 0 9292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_23
timestamp 1694700623
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1694700623
transform -1 0 9292 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_24
timestamp 1694700623
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1694700623
transform -1 0 9292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_25
timestamp 1694700623
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1694700623
transform -1 0 9292 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_26
timestamp 1694700623
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1694700623
transform -1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_27
timestamp 1694700623
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1694700623
transform -1 0 9292 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_28
timestamp 1694700623
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1694700623
transform -1 0 9292 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_29
timestamp 1694700623
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1694700623
transform -1 0 9292 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  rebuffer1
timestamp 1694700623
transform -1 0 4048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  rebuffer3
timestamp 1694700623
transform -1 0 4416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1694700623
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_31
timestamp 1694700623
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_32
timestamp 1694700623
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_33
timestamp 1694700623
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_34
timestamp 1694700623
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_35
timestamp 1694700623
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_36
timestamp 1694700623
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_37
timestamp 1694700623
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_38
timestamp 1694700623
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_39
timestamp 1694700623
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_40
timestamp 1694700623
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_41
timestamp 1694700623
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_42
timestamp 1694700623
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_43
timestamp 1694700623
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_44
timestamp 1694700623
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_45
timestamp 1694700623
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_46
timestamp 1694700623
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_47
timestamp 1694700623
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_48
timestamp 1694700623
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_49
timestamp 1694700623
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_50
timestamp 1694700623
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_51
timestamp 1694700623
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_52
timestamp 1694700623
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_53
timestamp 1694700623
transform 1 0 6256 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_54
timestamp 1694700623
transform 1 0 8832 0 1 9792
box -38 -48 130 592
<< labels >>
flabel metal4 s 2627 2128 2947 10384 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4674 2128 4994 10384 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 6721 2128 7041 10384 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 8768 2128 9088 10384 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3696 9340 4016 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 5736 9340 6056 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 7776 9340 8096 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 9816 9340 10136 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1967 2128 2287 10384 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4014 2128 4334 10384 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6061 2128 6381 10384 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 8108 2128 8428 10384 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3036 9340 3356 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 5076 9340 5396 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 7116 9340 7436 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 9156 9340 9476 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal2 s 5814 11802 5870 12602 0 FreeSans 224 90 0 0 clkout
port 3 nsew signal tristate
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 reset
port 4 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 sel[0]
port 5 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 sel[1]
port 6 nsew signal input
rlabel metal1 5198 9792 5198 9792 0 VGND
rlabel metal1 5198 10336 5198 10336 0 VPWR
rlabel metal1 7666 6358 7666 6358 0 _000_
rlabel metal1 6240 3094 6240 3094 0 _001_
rlabel via1 7677 6766 7677 6766 0 _002_
rlabel metal1 7079 2414 7079 2414 0 _003_
rlabel metal1 5520 9078 5520 9078 0 _004_
rlabel metal1 3450 2618 3450 2618 0 _005_
rlabel metal1 2157 5678 2157 5678 0 _006_
rlabel metal1 1748 6970 1748 6970 0 _007_
rlabel metal1 1472 8602 1472 8602 0 _008_
rlabel metal2 2898 9350 2898 9350 0 _009_
rlabel metal2 4370 9078 4370 9078 0 _010_
rlabel via1 7677 9622 7677 9622 0 _011_
rlabel metal1 7528 8534 7528 8534 0 _012_
rlabel metal1 1886 3706 1886 3706 0 _013_
rlabel metal1 1840 2618 1840 2618 0 _014_
rlabel via1 5754 3026 5754 3026 0 _015_
rlabel metal1 1656 8534 1656 8534 0 _016_
rlabel metal1 2714 7310 2714 7310 0 _017_
rlabel metal2 3174 9010 3174 9010 0 _018_
rlabel metal1 2990 8602 2990 8602 0 _019_
rlabel metal1 3174 7854 3174 7854 0 _020_
rlabel metal1 3772 8058 3772 8058 0 _021_
rlabel metal1 4876 8058 4876 8058 0 _022_
rlabel metal1 4094 8500 4094 8500 0 _023_
rlabel metal1 8004 9894 8004 9894 0 _024_
rlabel metal2 7498 9554 7498 9554 0 _025_
rlabel metal2 7222 8483 7222 8483 0 _026_
rlabel metal1 7866 10030 7866 10030 0 _027_
rlabel metal1 6900 9146 6900 9146 0 _028_
rlabel metal2 7314 9622 7314 9622 0 _029_
rlabel metal1 6946 8534 6946 8534 0 _030_
rlabel metal1 7590 8466 7590 8466 0 _031_
rlabel metal1 7774 3366 7774 3366 0 _032_
rlabel metal2 7314 8262 7314 8262 0 _033_
rlabel metal1 2346 3502 2346 3502 0 _034_
rlabel metal1 2346 3706 2346 3706 0 _035_
rlabel metal2 5382 4420 5382 4420 0 _036_
rlabel metal1 1978 3604 1978 3604 0 _037_
rlabel metal1 1610 2448 1610 2448 0 _038_
rlabel metal2 2346 3264 2346 3264 0 _039_
rlabel metal1 4002 2448 4002 2448 0 _040_
rlabel metal1 4416 3162 4416 3162 0 _041_
rlabel metal1 2162 2482 2162 2482 0 _042_
rlabel metal2 5474 2587 5474 2587 0 _043_
rlabel metal1 4186 2618 4186 2618 0 _044_
rlabel metal1 4554 3638 4554 3638 0 _045_
rlabel metal1 5750 2414 5750 2414 0 _046_
rlabel metal1 5152 5882 5152 5882 0 _047_
rlabel metal1 2438 7820 2438 7820 0 _048_
rlabel metal2 2714 8126 2714 8126 0 _049_
rlabel metal1 5244 10030 5244 10030 0 _050_
rlabel metal1 3542 5678 3542 5678 0 _051_
rlabel metal1 8602 5236 8602 5236 0 _052_
rlabel metal1 8648 5338 8648 5338 0 _053_
rlabel metal1 4922 4726 4922 4726 0 _054_
rlabel metal2 6854 4828 6854 4828 0 _055_
rlabel metal1 5750 7310 5750 7310 0 _056_
rlabel metal1 5842 7412 5842 7412 0 _057_
rlabel metal1 6578 6324 6578 6324 0 _058_
rlabel metal2 1702 9724 1702 9724 0 _059_
rlabel metal1 1702 7786 1702 7786 0 _060_
rlabel metal1 6118 6732 6118 6732 0 _061_
rlabel metal1 5658 6766 5658 6766 0 _062_
rlabel metal1 4554 5644 4554 5644 0 _063_
rlabel metal2 4554 6256 4554 6256 0 _064_
rlabel metal1 5198 3468 5198 3468 0 _065_
rlabel metal1 6808 5882 6808 5882 0 _066_
rlabel metal1 6302 4250 6302 4250 0 _067_
rlabel metal1 7866 3638 7866 3638 0 _068_
rlabel metal1 7820 3706 7820 3706 0 _069_
rlabel metal1 5658 4080 5658 4080 0 _070_
rlabel metal1 3542 7718 3542 7718 0 _071_
rlabel metal1 5198 9894 5198 9894 0 _072_
rlabel metal1 6486 6256 6486 6256 0 _073_
rlabel metal1 5750 2550 5750 2550 0 _074_
rlabel metal1 7682 7378 7682 7378 0 _075_
rlabel via2 7314 7395 7314 7395 0 _076_
rlabel metal1 7084 4590 7084 4590 0 _077_
rlabel metal1 7636 5746 7636 5746 0 _078_
rlabel metal1 7945 5610 7945 5610 0 _079_
rlabel metal2 7498 6018 7498 6018 0 _080_
rlabel metal1 7130 7276 7130 7276 0 _081_
rlabel metal1 7222 4624 7222 4624 0 _082_
rlabel metal1 7636 4250 7636 4250 0 _083_
rlabel metal1 6302 3536 6302 3536 0 _084_
rlabel metal2 7222 9792 7222 9792 0 _085_
rlabel metal1 5428 10166 5428 10166 0 _086_
rlabel metal1 5566 5882 5566 5882 0 _087_
rlabel metal2 5842 8653 5842 8653 0 _088_
rlabel metal1 3864 4794 3864 4794 0 _089_
rlabel metal1 5060 3502 5060 3502 0 _090_
rlabel metal1 4324 4454 4324 4454 0 _091_
rlabel metal2 5198 7106 5198 7106 0 _092_
rlabel metal2 7774 7905 7774 7905 0 _093_
rlabel metal1 5566 9010 5566 9010 0 _094_
rlabel metal1 2254 6426 2254 6426 0 _095_
rlabel metal2 3496 2516 3496 2516 0 _096_
rlabel metal1 3358 6222 3358 6222 0 _097_
rlabel metal1 3312 5338 3312 5338 0 _098_
rlabel viali 1641 6324 1641 6324 0 _099_
rlabel metal1 2990 6188 2990 6188 0 _100_
rlabel metal1 1886 6834 1886 6834 0 _101_
rlabel metal2 3542 6290 3542 6290 0 _102_
rlabel metal2 4462 7973 4462 7973 0 clk
rlabel metal1 5658 6426 5658 6426 0 clknet_0_clk
rlabel metal2 1426 5440 1426 5440 0 clknet_1_0__leaf_clk
rlabel metal2 1426 8160 1426 8160 0 clknet_1_1__leaf_clk
rlabel metal1 6164 10234 6164 10234 0 clkout
rlabel via1 3634 4998 3634 4998 0 cnt1\[0\]
rlabel metal1 3864 5202 3864 5202 0 cnt1\[1\]
rlabel metal1 1886 9690 1886 9690 0 cnt1\[2\]
rlabel metal1 1702 9418 1702 9418 0 cnt1\[3\]
rlabel metal1 3082 8364 3082 8364 0 cnt1\[4\]
rlabel metal1 2254 7888 2254 7888 0 cnt1\[5\]
rlabel metal1 8050 7888 8050 7888 0 cnt2\[0\]
rlabel metal2 7498 7735 7498 7735 0 cnt2\[1\]
rlabel metal1 2530 3536 2530 3536 0 cnt3\[0\]
rlabel metal2 3128 2516 3128 2516 0 cnt3\[1\]
rlabel metal1 4140 2550 4140 2550 0 cnt3\[2\]
rlabel metal1 8464 6426 8464 6426 0 cnt4\[0\]
rlabel metal1 7590 5338 7590 5338 0 cnt4\[1\]
rlabel metal2 8786 7140 8786 7140 0 cnt4\[2\]
rlabel metal1 8280 2958 8280 2958 0 cnt4\[3\]
rlabel metal1 5842 4624 5842 4624 0 net1
rlabel metal1 5336 2414 5336 2414 0 net13
rlabel metal2 2806 2587 2806 2587 0 net14
rlabel metal1 7038 8466 7038 8466 0 net15
rlabel metal1 3634 9894 3634 9894 0 net16
rlabel metal1 2530 2448 2530 2448 0 net17
rlabel metal1 2622 4556 2622 4556 0 net2
rlabel metal1 7682 3162 7682 3162 0 net20
rlabel metal2 7038 3910 7038 3910 0 net21
rlabel metal1 8280 7514 8280 7514 0 net22
rlabel metal1 2047 8466 2047 8466 0 net23
rlabel metal1 7406 6766 7406 6766 0 net24
rlabel metal1 2530 4624 2530 4624 0 net3
rlabel metal1 6486 9962 6486 9962 0 net4
rlabel metal2 1610 7378 1610 7378 0 net5
rlabel metal2 3358 7140 3358 7140 0 net6
rlabel metal2 4370 6426 4370 6426 0 net7
rlabel metal2 5658 9146 5658 9146 0 net9
rlabel metal3 1004 6188 1004 6188 0 reset
rlabel metal1 1932 2414 1932 2414 0 sel[0]
rlabel metal2 5198 1554 5198 1554 0 sel[1]
<< properties >>
string FIXED_BBOX 0 0 10458 12602
<< end >>
